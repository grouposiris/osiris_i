// This is the unpowered netlist.
module core (clk,
    o_mem_write_M,
    rst,
    i_instr_ID,
    i_read_data_M,
    o_data_addr_M,
    o_funct3_MEM,
    o_pc_IF,
    o_write_data_M);
 input clk;
 output o_mem_write_M;
 input rst;
 input [31:0] i_instr_ID;
 input [31:0] i_read_data_M;
 output [31:0] o_data_addr_M;
 output [2:0] o_funct3_MEM;
 output [31:0] o_pc_IF;
 output [31:0] o_write_data_M;

 wire net476;
 wire net477;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ;
 wire \U_CONTROL_UNIT.i_branch_EX ;
 wire \U_CONTROL_UNIT.i_jump_EX ;
 wire \U_DATAPATH.U_EX_MEM.i_funct3_EX[0] ;
 wire \U_DATAPATH.U_EX_MEM.i_funct3_EX[1] ;
 wire \U_DATAPATH.U_EX_MEM.i_funct3_EX[2] ;
 wire \U_DATAPATH.U_EX_MEM.i_mem_write_EX ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[10] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[11] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[12] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[13] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[14] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[15] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[16] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[17] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[18] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[19] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[20] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[21] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[22] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[23] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[24] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[25] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[26] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[27] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[28] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[29] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[2] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[30] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[31] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[3] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[4] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[5] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[6] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[7] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[8] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[9] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[0] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[1] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[2] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[3] ;
 wire \U_DATAPATH.U_EX_MEM.i_reg_write_EX ;
 wire \U_DATAPATH.U_EX_MEM.i_result_src_EX[0] ;
 wire \U_DATAPATH.U_EX_MEM.i_result_src_EX[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[10] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[11] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[12] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[13] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[14] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[15] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[16] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[17] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[18] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[19] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[20] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[21] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[22] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[23] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[24] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[25] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[26] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[27] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[28] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[29] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[30] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[31] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[4] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[5] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[6] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[7] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[8] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[9] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[10] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[11] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[12] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[13] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[14] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[15] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[16] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[17] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[18] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[19] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[20] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[21] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[22] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[23] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[24] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[25] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[26] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[27] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[28] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[29] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[30] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[31] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[4] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[5] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[6] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[7] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[8] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[9] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_reg_write_M ;
 wire \U_DATAPATH.U_EX_MEM.o_result_src_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_result_src_M[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[0] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[1] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[0] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[1] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[0] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[1] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.o_addr_src_EX ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_src_EX ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[9] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[9] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[9] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[10] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[11] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[12] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[13] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[14] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[15] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[16] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[17] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[18] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[19] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[20] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[21] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[22] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[23] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[24] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[25] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[26] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[27] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[28] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[29] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[2] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[30] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[31] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[3] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[4] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[5] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[6] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[7] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[8] ;
 wire \U_DATAPATH.U_IF_ID.i_pc_IF[9] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[10] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[11] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[12] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[13] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[14] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[15] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[16] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[17] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[18] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[19] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[20] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[21] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[22] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[23] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[24] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[25] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[26] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[27] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[28] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[29] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[2] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[30] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[31] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[3] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[4] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[5] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[6] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[7] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[8] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[9] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[11] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[19] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[24] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[25] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[26] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[27] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[28] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[29] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[1] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[1] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_9_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net21;
 wire net210;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net211;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net212;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net213;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net216;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net217;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net218;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net219;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net22;
 wire net220;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net221;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net222;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net223;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net235;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net236;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net237;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net238;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net239;
 wire net2390;
 wire net2391;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\U_DATAPATH.U_ID_EX.i_rs2_ID[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\U_DATAPATH.U_ID_EX.o_pc_EX[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_1596_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\U_DATAPATH.U_ID_EX.o_pc_EX[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net2251));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\U_DATAPATH.U_ID_EX.o_pc_EX[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__B (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__B (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__B (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__B (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__S0 (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__S1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A2 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__B1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__B (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A2 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__B1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__A_N (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__A_N (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__B (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__B1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__B2 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A1 (.DIODE(net1996));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__A (.DIODE(net1996));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__B1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__B (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__B (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__B (.DIODE(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__C (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__A1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__B1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A1 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__B1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__B (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__B (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__A_N (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__B1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__B2 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A2 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__B1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__B (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__B (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__B2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__B (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__A1 (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A1 (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__B (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__B1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__B1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__B (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__B (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__B (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__B1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__B (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__B (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A_N (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__C (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__B1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__B1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__B (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__B (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__B (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A_N (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__C (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__B1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__B1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A_N (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__C (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A1 (.DIODE(net2185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__B1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A1 (.DIODE(_1444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__B1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A_N (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__B2 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A2 (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A_N (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__C (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__B1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__B1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__A_N (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__B1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__B2 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A1 (.DIODE(net2006));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A2 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A (.DIODE(net2006));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__B1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__B (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__B (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A_N (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__C (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__B1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A1 (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__B1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__B (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__B (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__A_N (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__B1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__B2 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__A1 (.DIODE(net2159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A2 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__B1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__A_N (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__B1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__B2 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A1 (.DIODE(net2178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__A (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__B1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__B (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__B (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__C (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A1 (.DIODE(net1984));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__B1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A2 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A2 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__B (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__B (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A_N (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__C (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__B1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A2 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__A2 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__B (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__B (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__B (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A2 (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__C (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__B (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__C (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A3 (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__B1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A1 (.DIODE(net2350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__B1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__B (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__B (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__A2 (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__C (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__B1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__A1 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__A (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__B (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__B (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__A_N (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A1 (.DIODE(net2034));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__B1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A0 (.DIODE(net2160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A1 (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__B1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__A (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__B (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__B (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__C (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A1 (.DIODE(net1928));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__B1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__B (.DIODE(net2229));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A2 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A2 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A (.DIODE(net1928));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__B1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__B (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__B (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A1 (.DIODE(net2067));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__B1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A1 (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__B1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__B (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__B (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__B (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__A1 (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A1 (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__B (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__C (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__C (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__B1 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__B (.DIODE(net2170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A (.DIODE(_1612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__B1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__A (.DIODE(_1612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__C (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__A1 (.DIODE(_1612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__B1 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__B (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__C (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A1 (.DIODE(net2104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__B1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A1 (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__B1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__B (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__B (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__C (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__B1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A1 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__B (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__C (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A2 (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__B1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__B2 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__A (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__B (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__B (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__B (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__B2 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A1 (.DIODE(net2008));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__B (.DIODE(net2224));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__A2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__B (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__C (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__B (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__B (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__C (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__A1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__B1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__A0 (.DIODE(net2214));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__A1 (.DIODE(_1657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__B (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__A (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__B (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__C (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__B1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__A1 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__B1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__B (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__B (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__B (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__B1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__A1 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A2 (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__B2 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__B (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__B (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A_N (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__B1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__B2 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__A2 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__B1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__B (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__B (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__A_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__B (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__C (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__B1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__A1 (.DIODE(_1704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__B (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__C (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__B1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__B (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__B (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A_N (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__B (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A_N (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__B1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__C1 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__A_N (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__B (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__B (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A_N (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__B (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__A_N (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__B (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__B (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A_N (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__B (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__A_N (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A3 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__B1 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A_N (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A_N (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__A2 (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__B1 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__A_N (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__B (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A_N (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__C1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__A_N (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__B1 (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A_N (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__B1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A2 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A3 (.DIODE(_1765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A0 (.DIODE(\U_DATAPATH.U_ID_EX.o_pc_EX[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__B (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__C (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__A2 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__B (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__C (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__A (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__A (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__B (.DIODE(_1795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__A1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__A2 (.DIODE(_1795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__S (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__A (.DIODE(_1795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A0 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__S (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__B (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__A (.DIODE(net2229));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__A (.DIODE(net2229));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__S (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A (.DIODE(net2170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A (.DIODE(net2170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__S (.DIODE(\U_DATAPATH.U_ID_EX.o_addr_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__A (.DIODE(net2160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__A (.DIODE(net2160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__S (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__A (.DIODE(net2224));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__S (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__A0 (.DIODE(_1858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__S (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__S (.DIODE(\U_DATAPATH.U_ID_EX.o_addr_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__S (.DIODE(\U_DATAPATH.U_ID_EX.o_addr_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__A (.DIODE(net2214));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__S (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__A0 (.DIODE(_1885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__S (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__S (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__B (.DIODE(_1886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__S (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__S (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__B (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__S (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__B (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__B (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A0 (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__B (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__A_N (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__S (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__A0 (.DIODE(\U_DATAPATH.U_ID_EX.o_pc_EX[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__A2 (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__B (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__C (.DIODE(_1959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__S (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__S (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__S (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__C (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__S (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__S (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__S (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__S (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__S (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__S (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__S (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__S (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__B (.DIODE(_2074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__B (.DIODE(_2074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__A1 (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__B1 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__B1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__A2 (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__B1 (.DIODE(_1959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__B1 (.DIODE(_2099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__B (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__S (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__B (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__A3 (.DIODE(_1886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__B (.DIODE(_1886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__S (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__S (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__A2 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__B (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__S (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__S (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__S (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__S (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__S (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__A1 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__S (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__S (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__S (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__A1 (.DIODE(_1959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__S (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__A1 (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__S (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__S (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__A1 (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__S (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__S (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__S (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__A1 (.DIODE(_1886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__S (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__S (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__S (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__S (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__S (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__S (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__S (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__S (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__A1 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__S (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__S (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__S (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__S (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__S (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__S (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__S (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__S (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__S (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__S (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__S (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__S (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__S0 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__S0 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__S0 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__S0 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__S (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__S (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__S (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__S (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__S (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__S (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__S (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__S (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__S (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__S (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__S1 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__S (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__S (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__S1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__S (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__S (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__S1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__S (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__S1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__S1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__S1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__S1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__S1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__S1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__S1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__S1 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__S1 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__S1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__S0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__S1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__S0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__S (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__C_N (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__B (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__B (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__S (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__C_N (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__S (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__C_N (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A (.DIODE(net2151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A (.DIODE(net2153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A (.DIODE(net2107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A (.DIODE(net1998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A (.DIODE(net1990));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A (.DIODE(net2126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__B (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__B1 (.DIODE(_2522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__B1 (.DIODE(_2522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A (.DIODE(net2018));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A (.DIODE(net1972));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A (.DIODE(net2116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A (.DIODE(net1742));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A (.DIODE(net2073));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__A (.DIODE(net1945));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__B (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__B (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A2 (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A2 (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__B1 (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A (.DIODE(net1990));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__B (.DIODE(net1998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__C (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__A_N (.DIODE(net1990));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A (.DIODE(net1998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__B (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__B (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__B (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A (.DIODE(net1990));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A (.DIODE(net1990));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A (.DIODE(net1998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__B (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__B (.DIODE(net2197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__C_N (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A1 (.DIODE(net1990));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A2 (.DIODE(net1998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A (.DIODE(net1998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__B (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A1 (.DIODE(net1998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A2 (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A (.DIODE(net1990));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__B (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__B (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__C (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__C (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__C (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__C (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__C (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__C (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__C (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__C (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__C (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__C (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__C (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__C (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__C (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__C (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__C (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__C (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__C (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__C (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__C (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__C (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__C (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__C (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__C (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__C (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__C (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__C (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__C (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__C (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__C (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__C (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__C (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__C (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__A (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__C (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__C (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__C (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__C (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__C (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__B (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__C (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__C (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__C (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__C (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__C (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__B (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__C (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__B (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__B (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__B (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__B (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__B (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__C (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__C (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__B (.DIODE(net2122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__B (.DIODE(net2122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__C (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__C (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__C (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__C (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__C (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__C (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A (.DIODE(\U_DATAPATH.U_ID_EX.i_rs1_ID[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__C (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__C (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__C (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__C (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__B (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__C (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__B (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__B (.DIODE(net2122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__C (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__C (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__C (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__C (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A (.DIODE(\U_DATAPATH.U_ID_EX.i_rs1_ID[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A (.DIODE(net2151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A (.DIODE(net2153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__C (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A (.DIODE(net2107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__C (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A2 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__B (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__B (.DIODE(_1858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__B (.DIODE(_1885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__B (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__B (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__B (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__B (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__B (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A0 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A1 (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A2 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A3 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A0 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A1 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A2 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A3 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__S0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A0 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A1 (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A0 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A1 (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A3 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__A0 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__A1 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__A0 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__A1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__S (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A0 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A0 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__A1 (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A0 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A0 (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A1 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A0 (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__S (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__C (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__D (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__B1 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__B1 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__A (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__C (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__B (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__C (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__B2 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__C1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A0 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A0 (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A0 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A1 (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__B (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A1 (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__A2 (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A1 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__B2 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__C (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__B1 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__B1 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A0 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A1 (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__S (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__B1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__B2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__C1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A0 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A1 (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A1_N (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__B2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A0 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A1 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A2 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A3 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__S1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A0 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A1 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A3 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__S1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A0 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A1 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A0 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A0 (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A1 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A0 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A1 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A2 (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A3 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__S0 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__S (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A2 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A0 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A1 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__S (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A0 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A1 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A2 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A3 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__S0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A0 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A1 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A2 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A3 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__S0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__B2 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__B (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__B1 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A2 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__C1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A1 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__B2 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__B (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__A (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A0 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A1 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__B1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__C1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__B2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A0 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A1 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A2 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A3 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A0 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A3 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__S0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__S (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__A2 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__B (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A2 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__B1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__A0 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__A1 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__A2 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__A3 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__C1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__C1 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__B1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__C1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A0 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A1 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__S (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__B2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__B1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A1 (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__B1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__A1 (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A1 (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A2 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5913__A (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A0 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A1 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A2 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A3 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__B (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__B (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__C1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__C (.DIODE(_2947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__C1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__B (.DIODE(_2953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A0 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A1 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__A1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__A2 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__B1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A1_N (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__A1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__C1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A2 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__C1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A2 (.DIODE(_2953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A0 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A1 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A2 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A3 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__S (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A1 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__B2 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__B1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__C1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__C1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A1 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__A (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A0 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A1 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__S (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__A1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__B2 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__A1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__B1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__A1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__A1_N (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__B2 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__A1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6004__C1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__A (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__A (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A0 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A1 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A3 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__S0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__A (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__A1 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__B1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__C1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__A1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__C1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__C1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6026__A (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6026__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__A (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__A (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A0 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A1 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A2 (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A3 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A2 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__B2 (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__C1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__A1_N (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__A1 (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__A2 (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__A (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__A (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A1 (.DIODE(_3059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__B1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__A1 (.DIODE(_3059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A0 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A1 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A3 (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__B2 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A1_N (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__B1 (.DIODE(_3076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__C1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__C1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__A (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__A (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__A1 (.DIODE(_3059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__B1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A0 (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A1 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A2 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A3 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__B1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__C1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__B2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A1_N (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A2 (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A2 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__B1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__C1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__A (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__B1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A0 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A1 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A2 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A3 (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__S0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__A1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A2 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__A2 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__B2 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__A2 (.DIODE(_3113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__C1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__B1 (.DIODE(_3117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__B2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__C1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__A (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A0 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A1 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A2 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A3 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__B1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__C1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__B1 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__B2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__B1 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__A1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__B1 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__B1 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A1 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__C1 (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A2 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__B1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__B (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__A (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__A (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A0 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A1 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A2 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A3 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__S0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__B (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__A2 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__B1 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__A2 (.DIODE(_3152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__D1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A2 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A3 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__S1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__S (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__B1 (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__C1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__A2 (.DIODE(_3152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__B2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__B2 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__C1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__B1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__B1 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__B2 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__C1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A0 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A2 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__A1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A1 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__B2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__B1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A1 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__A (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__A (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A2 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A3 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__S (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__B1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__B2 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__C1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__A2 (.DIODE(_3152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__B2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__A1 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__B2 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__A1 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__A2 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__B1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__C1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A2 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__S0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__B1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__B1 (.DIODE(_3152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__B1 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__B1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__B1 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__A2 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__C1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A0 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6236__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__C1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__B1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__C1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__B1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__A3 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__S0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__A1_N (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__B1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__C1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6258__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__D1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__C1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__A2 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__C1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__B2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A1 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__C1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6280__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__B1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A1_N (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__B1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__C1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__B1 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__A2 (.DIODE(_3152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__C1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__A (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__A (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__A1 (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__C1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A2 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__C1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__B2 (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__B2 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__A2 (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__C1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6318__A (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__A (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A0 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A2 (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__S (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__B2 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__A1_N (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__B2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A2 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__B1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__C1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__A (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__A (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__B1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__A0 (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__A2 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__A3 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__A1_N (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__B1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A2 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__C1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__B2 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__C1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__A (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__A (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A0 (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A2 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A3 (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__B1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__C1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__C1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__A (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A0 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A2 (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A3 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__A1_N (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A2 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__C1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__B2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A2 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__C1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__B (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__A (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A0 (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A1 (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A2 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A3 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__S1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__S (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__B2 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__B1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__C1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__A2 (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__D1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__C1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__C1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A0 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A1 (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A2 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A3 (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__S1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__C1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A2 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__C1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__A2 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__B1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__A1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__A2 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__C1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__A3 (.DIODE(_3152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A2 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__C1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__B (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__A3 (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__B1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__B (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__B (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__B1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__B (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__B (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__B (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__B (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__B (.DIODE(_1657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__B (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__B (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__B (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__B (.DIODE(_1704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__B1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__B (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__B (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__B (.DIODE(_1444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__B (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__B (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__B (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__B (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__B (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__B (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__B (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__B (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__S (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__6461__S (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__S (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__S (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6505__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__B (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__B (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__A (.DIODE(net1984));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__A (.DIODE(net1928));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__A (.DIODE(net2067));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__B (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__A (.DIODE(net2034));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__A (.DIODE(net2008));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__A (.DIODE(net2104));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__B (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__B (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__B (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__B (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__B (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6544__B (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__B (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__A (.DIODE(net2185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__B (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__A (.DIODE(net2159));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__B (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__A (.DIODE(net2006));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__A (.DIODE(net2178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__B (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__A (.DIODE(net1996));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__B (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__A (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__B (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__A (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__A (.DIODE(net1998));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__C (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__A (.DIODE(net1990));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__C (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__C (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A3 (.DIODE(_3418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__A (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__B (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A3 (.DIODE(_3418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A1 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__A1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__C (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A1 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__A (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__A3 (.DIODE(_3461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A3 (.DIODE(_3461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__A1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__A1 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__B (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6842__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6845__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6846__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6846__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6846__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6862__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6862__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__C (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6881__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6881__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__A3 (.DIODE(_3503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__A1 (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__A3 (.DIODE(_3503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__A1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__A1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__A1 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6924__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6926__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__A (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__C (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__A1 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__A2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__A (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__A (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6948__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6948__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__A3 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__A (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__A1 (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__A (.DIODE(_1596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6958__A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6958__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__A (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__6962__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__A (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6964__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6964__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__A (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__A (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6968__A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6968__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__A (.DIODE(_1702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__6976__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6976__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6978__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6978__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6981__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__6982__A1 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6982__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__6984__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6984__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__A (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6988__A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6988__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__6990__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__A (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__6992__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__A (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__6998__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6998__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__A (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__A (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__A (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__A (.DIODE(net1990));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__B (.DIODE(net1998));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__C (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__A1_N (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__A1 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__C1 (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__A1 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__A2 (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__C1 (.DIODE(net1998));
 sky130_fd_sc_hd__diode_2 ANTENNA__7018__A (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7019__A1 (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7019__B2 (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7023__A1 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__A0 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__A (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__A1 (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__B2 (.DIODE(net2205));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__A0 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__7033__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__7041__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__7048__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__7054__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__7059__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__7061__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__7065__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__A (.DIODE(net1945));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__B (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__C (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__A (.DIODE(net1945));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__A (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__B (.DIODE(net2001));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__A1 (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__A (.DIODE(net2073));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__B (.DIODE(net2001));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__A1 (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7072__A (.DIODE(net1742));
 sky130_fd_sc_hd__diode_2 ANTENNA__7072__B (.DIODE(net2001));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__A1 (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7074__A (.DIODE(net2116));
 sky130_fd_sc_hd__diode_2 ANTENNA__7074__B (.DIODE(net2001));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__A1 (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__A2 (.DIODE(_3596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__A (.DIODE(net1972));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__B (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__A1 (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__A (.DIODE(net2018));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__B (.DIODE(net2001));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__A1 (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__A (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__B (.DIODE(net2001));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__A1 (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7082__A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__7082__B (.DIODE(net2001));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__A1 (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__A (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__B (.DIODE(net2001));
 sky130_fd_sc_hd__diode_2 ANTENNA__7085__A1 (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7085__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__B (.DIODE(net2001));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__A1 (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__B (.DIODE(net2001));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__A1 (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__A (.DIODE(net2126));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__A (.DIODE(net1945));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7093__A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__7098__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__A (.DIODE(net1990));
 sky130_fd_sc_hd__diode_2 ANTENNA__7102__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__A (.DIODE(net1998));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7105__A (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__A1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__B2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA__7109__B1 (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__A (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__C (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__A (.DIODE(net2073));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__C (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__A (.DIODE(net1742));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__C (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__A (.DIODE(net2116));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__C (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__A (.DIODE(net1972));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__C (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__A (.DIODE(net2018));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__C (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__A1 (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7118__B2 (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__7119__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__7119__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7120__A1 (.DIODE(net2107));
 sky130_fd_sc_hd__diode_2 ANTENNA__7120__B2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__7121__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__7121__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__A1 (.DIODE(net2153));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__B2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__A1 (.DIODE(net2151));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__B2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__A1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__B2 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7133__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7136__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7137__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7139__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7140__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7146__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7147__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7148__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7149__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7150__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7152__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__7159__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__7225__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7227__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7229__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7230__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7231__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__7232__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7233__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7234__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7235__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7236__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7239__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7240__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7241__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7242__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__7247__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7249__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7250__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7251__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7260__CLK (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7286__RESET_B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__7634__D (.DIODE(_0511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7705__D (.DIODE(_0582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7734__D (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7757__D (.DIODE(_0634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7762__D (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7840__D (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7845__D (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7850__D (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7855__D (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7858__D (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7876__D (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7877__D (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7879__D (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7884__CLK (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7884__D (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7891__D (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7893__D (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7894__D (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7897__D (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7898__D (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7902__D (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7905__D (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7976__D (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__8010__D (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8041__D (.DIODE(_0052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8402__D (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8421__D (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(_2522_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(_2522_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(_2522_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(_3500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(_3500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(_3458_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(_3458_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(_3453_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(_3453_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(_2644_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(_2644_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(_2635_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(_2635_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(_2620_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(_2620_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(_3503_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(_3498_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(_3498_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(_3496_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(_3496_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(_3461_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(_3461_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(_3451_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(_3451_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_A (.DIODE(_2075_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(_2075_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_A (.DIODE(_3494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(_3494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(_3418_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout311_A (.DIODE(_3418_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout312_A (.DIODE(_3417_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout313_A (.DIODE(_3417_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout314_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout317_A (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout318_A (.DIODE(_1702_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout319_A (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout322_A (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout324_A (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout325_A (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout326_A (.DIODE(_1596_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout327_A (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout331_A (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout332_A (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout333_A (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout334_A (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout335_A (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout339_A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout340_A (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout345_A (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout346_A (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout347_A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout348_A (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout351_A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout353_A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout360_A (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout361_A (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout364_A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout365_A (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout366_A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout368_A (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout369_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout371_A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout373_A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout375_A (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout376_A (.DIODE(\U_DATAPATH.U_ID_EX.o_addr_src_EX ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout379_A (.DIODE(net2112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout380_A (.DIODE(net2112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout381_A (.DIODE(net2098));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout382_A (.DIODE(net2098));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout383_A (.DIODE(net2098));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout384_A (.DIODE(net2098));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout385_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout386_A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout387_A (.DIODE(net2096));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout388_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout389_A (.DIODE(net2096));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout390_A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout391_A (.DIODE(net2096));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout392_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout393_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout394_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout395_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout396_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout397_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout398_A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout399_A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout401_A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout402_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout403_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout404_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout405_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout407_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout408_A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout410_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout411_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout412_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout413_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout415_A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout416_A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout417_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout418_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout419_A (.DIODE(net2174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout420_A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout421_A (.DIODE(net2174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout422_A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout423_A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout424_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout425_A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout426_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout427_A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout428_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout429_A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout430_A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout431_A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout432_A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout433_A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout435_A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout436_A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout437_A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout438_A (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout439_A (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout440_A (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout441_A (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout442_A (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout443_A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout444_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout445_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout446_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout447_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout448_A (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout449_A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout450_A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout451_A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout452_A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout453_A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout454_A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout455_A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout456_A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout457_A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout458_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout459_A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout460_A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout461_A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout462_A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout463_A (.DIODE(_0069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout464_A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout465_A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout466_A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout467_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout468_A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout469_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout470_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout471_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout472_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold100_A (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1155_A (.DIODE(net2205));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1170_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1237_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1254_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1307_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1358_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1400_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1401_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1417_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1434_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1452_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1454_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1455_A (.DIODE(net2197));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1468_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1469_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1483_A (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1490_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1492_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1503_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1515_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1523_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1526_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1541_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1542_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1545_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1552_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1553_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1555_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1563_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1567_A (.DIODE(\U_DATAPATH.U_IF_ID.o_instr_ID[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1569_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1574_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1576_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1577_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1579_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1580_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1582_A (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1609_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1615_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1616_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1625_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1631_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1635_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1636_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1642_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1654_A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1655_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1662_A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1672_A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1678_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1679_A (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1681_A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1689_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1699_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1708_A (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1755_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1757_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1786_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1788_A (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1793_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1802_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1803_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1807_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1808_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1810_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1812_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1814_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1816_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1817_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1820_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1821_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1822_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1827_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1828_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1829_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1830_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1831_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1832_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1834_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1835_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1839_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1840_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1844_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1847_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold355_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold874_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap355_A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire301_A (.DIODE(_2075_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_223_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_224_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _3632_ (.A(net2124),
    .Y(_1277_));
 sky130_fd_sc_hd__inv_2 _3633_ (.A(net2000),
    .Y(_1278_));
 sky130_fd_sc_hd__inv_2 _3634_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .Y(_1279_));
 sky130_fd_sc_hd__inv_2 _3635_ (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ),
    .Y(_1280_));
 sky130_fd_sc_hd__inv_2 _3636_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .Y(_1281_));
 sky130_fd_sc_hd__inv_2 _3637_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .Y(_1282_));
 sky130_fd_sc_hd__inv_2 _3638_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .Y(_1283_));
 sky130_fd_sc_hd__inv_2 _3639_ (.A(net378),
    .Y(_1284_));
 sky130_fd_sc_hd__inv_2 _3640_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .Y(_1285_));
 sky130_fd_sc_hd__inv_2 _3641_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ),
    .Y(_1286_));
 sky130_fd_sc_hd__inv_2 _3642_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ),
    .Y(_1287_));
 sky130_fd_sc_hd__inv_2 _3643_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ),
    .Y(_1288_));
 sky130_fd_sc_hd__inv_2 _3644_ (.A(net2075),
    .Y(_1289_));
 sky130_fd_sc_hd__inv_2 _3645_ (.A(net2066),
    .Y(_1290_));
 sky130_fd_sc_hd__inv_4 _3646_ (.A(net471),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _3647__1 (.A(clknet_leaf_38_clk),
    .Y(net480));
 sky130_fd_sc_hd__nand2b_1 _3648_ (.A_N(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .Y(_1291_));
 sky130_fd_sc_hd__and2b_1 _3649_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .B(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .X(_1292_));
 sky130_fd_sc_hd__nand2b_1 _3650_ (.A_N(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .Y(_1293_));
 sky130_fd_sc_hd__nor4_1 _3651_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .C(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .D(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .Y(_1294_));
 sky130_fd_sc_hd__a221o_1 _3652_ (.A1(_1279_),
    .A2(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .B1(_1280_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .C1(_1292_),
    .X(_1295_));
 sky130_fd_sc_hd__nand2_1 _3653_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .Y(_1296_));
 sky130_fd_sc_hd__or2_1 _3654_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .X(_1297_));
 sky130_fd_sc_hd__a21o_1 _3655_ (.A1(_1296_),
    .A2(_1297_),
    .B1(_1294_),
    .X(_1298_));
 sky130_fd_sc_hd__o2111ai_4 _3656_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .A2(_1280_),
    .B1(_1291_),
    .C1(_1293_),
    .D1(net2109),
    .Y(_1299_));
 sky130_fd_sc_hd__nor3_4 _3657_ (.A(_1295_),
    .B(_1298_),
    .C(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__or3_1 _3658_ (.A(_1295_),
    .B(_1298_),
    .C(_1299_),
    .X(_1301_));
 sky130_fd_sc_hd__nand2b_1 _3659_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .Y(_1302_));
 sky130_fd_sc_hd__and2b_1 _3660_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .X(_1303_));
 sky130_fd_sc_hd__nand2b_1 _3661_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .Y(_1304_));
 sky130_fd_sc_hd__nand2_1 _3662_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .Y(_1305_));
 sky130_fd_sc_hd__or2_1 _3663_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .X(_1306_));
 sky130_fd_sc_hd__a21o_1 _3664_ (.A1(_1305_),
    .A2(_1306_),
    .B1(_1294_),
    .X(_1307_));
 sky130_fd_sc_hd__a221o_1 _3665_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .A2(_1281_),
    .B1(_1283_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .C1(_1303_),
    .X(_1308_));
 sky130_fd_sc_hd__o2111a_1 _3666_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .A2(_1281_),
    .B1(_1302_),
    .C1(_1304_),
    .D1(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .X(_1309_));
 sky130_fd_sc_hd__nor3b_1 _3667_ (.A(_1307_),
    .B(_1308_),
    .C_N(_1309_),
    .Y(_1310_));
 sky130_fd_sc_hd__or3b_4 _3668_ (.A(_1307_),
    .B(_1308_),
    .C_N(_1309_),
    .X(_1311_));
 sky130_fd_sc_hd__nor2_8 _3669_ (.A(net355),
    .B(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__nor2_8 _3670_ (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(net435),
    .Y(_1313_));
 sky130_fd_sc_hd__or2_1 _3671_ (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(net436),
    .X(_1314_));
 sky130_fd_sc_hd__and2_1 _3672_ (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(net436),
    .X(_1315_));
 sky130_fd_sc_hd__mux4_2 _3673_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[31] ),
    .A1(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[31] ),
    .A2(net55),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[31] ),
    .S0(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .S1(net436),
    .X(_1316_));
 sky130_fd_sc_hd__nor2_1 _3674_ (.A(net354),
    .B(net349),
    .Y(_1317_));
 sky130_fd_sc_hd__a22o_1 _3675_ (.A1(_1312_),
    .A2(net368),
    .B1(net307),
    .B2(net2180),
    .X(_1318_));
 sky130_fd_sc_hd__a21oi_4 _3676_ (.A1(net2158),
    .A2(net354),
    .B1(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__nand2_1 _3677_ (.A(net2267),
    .B(net377),
    .Y(_1320_));
 sky130_fd_sc_hd__o21ai_4 _3678_ (.A1(net377),
    .A2(_1319_),
    .B1(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__or4_1 _3679_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ),
    .C(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ),
    .D(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ),
    .X(_1322_));
 sky130_fd_sc_hd__o2bb2a_2 _3680_ (.A1_N(_1288_),
    .A2_N(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .B1(_1280_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .X(_1323_));
 sky130_fd_sc_hd__o22a_1 _3681_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .A2(_1287_),
    .B1(_1288_),
    .B2(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .X(_1324_));
 sky130_fd_sc_hd__a22oi_1 _3682_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .A2(_1286_),
    .B1(_1287_),
    .B2(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .Y(_1325_));
 sky130_fd_sc_hd__o211a_1 _3683_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .A2(_1286_),
    .B1(_1322_),
    .C1(\U_DATAPATH.U_EX_MEM.o_reg_write_M ),
    .X(_1326_));
 sky130_fd_sc_hd__o2111a_2 _3684_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ),
    .A2(_1285_),
    .B1(_1324_),
    .C1(_1325_),
    .D1(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__and2b_1 _3685_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .X(_1328_));
 sky130_fd_sc_hd__a221o_1 _3686_ (.A1(_1281_),
    .A2(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ),
    .B1(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ),
    .B2(_1283_),
    .C1(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__xor2_1 _3687_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ),
    .X(_1330_));
 sky130_fd_sc_hd__a221o_1 _3688_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .A2(_1286_),
    .B1(_1288_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .C1(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__o211a_1 _3689_ (.A1(_1282_),
    .A2(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .B1(_1322_),
    .C1(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .X(_1332_));
 sky130_fd_sc_hd__or3b_2 _3690_ (.A(_1329_),
    .B(_1331_),
    .C_N(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__a21oi_4 _3691_ (.A1(net364),
    .A2(net347),
    .B1(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__and3_1 _3692_ (.A(net88),
    .B(net365),
    .C(net348),
    .X(_1335_));
 sky130_fd_sc_hd__a21boi_4 _3693_ (.A1(net364),
    .A2(net347),
    .B1_N(_1333_),
    .Y(_1336_));
 sky130_fd_sc_hd__a221o_4 _3694_ (.A1(net368),
    .A2(net305),
    .B1(net303),
    .B2(net2277),
    .C1(_1335_),
    .X(_1337_));
 sky130_fd_sc_hd__clkinv_4 _3695_ (.A(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__xnor2_4 _3696_ (.A(_1321_),
    .B(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__and2b_1 _3697_ (.A_N(net436),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[28] ),
    .X(_1340_));
 sky130_fd_sc_hd__and2b_1 _3698_ (.A_N(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(net436),
    .X(_1341_));
 sky130_fd_sc_hd__a221o_1 _3699_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[28] ),
    .A2(net370),
    .B1(net367),
    .B2(net51),
    .C1(_1340_),
    .X(_1342_));
 sky130_fd_sc_hd__mux2_2 _3700_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[28] ),
    .A1(_1342_),
    .S(net372),
    .X(_1343_));
 sky130_fd_sc_hd__a22o_1 _3701_ (.A1(net2274),
    .A2(net307),
    .B1(net346),
    .B2(_1312_),
    .X(_1344_));
 sky130_fd_sc_hd__a21oi_4 _3702_ (.A1(net1996),
    .A2(net354),
    .B1(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__nand2_1 _3703_ (.A(net377),
    .B(net2040),
    .Y(_1346_));
 sky130_fd_sc_hd__o21ai_4 _3704_ (.A1(net377),
    .A2(_1345_),
    .B1(_1346_),
    .Y(_1347_));
 sky130_fd_sc_hd__inv_2 _3705_ (.A(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__and3_1 _3706_ (.A(net1996),
    .B(net365),
    .C(net348),
    .X(_1349_));
 sky130_fd_sc_hd__a221o_4 _3707_ (.A1(net2270),
    .A2(net303),
    .B1(net346),
    .B2(net305),
    .C1(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__nand2_1 _3708_ (.A(_1347_),
    .B(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__or2_1 _3709_ (.A(_1347_),
    .B(_1350_),
    .X(_1352_));
 sky130_fd_sc_hd__and2b_1 _3710_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ),
    .X(_1353_));
 sky130_fd_sc_hd__a221o_1 _3711_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[30] ),
    .A2(net369),
    .B1(net366),
    .B2(net54),
    .C1(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__mux2_4 _3712_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[30] ),
    .A1(_1354_),
    .S(net371),
    .X(_1355_));
 sky130_fd_sc_hd__and3_1 _3713_ (.A(net351),
    .B(net349),
    .C(net345),
    .X(_1356_));
 sky130_fd_sc_hd__a221o_4 _3714_ (.A1(net670),
    .A2(net353),
    .B1(net306),
    .B2(net2312),
    .C1(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__mux2_2 _3715_ (.A0(net2313),
    .A1(_1357_),
    .S(net374),
    .X(_1358_));
 sky130_fd_sc_hd__and3_1 _3716_ (.A(net87),
    .B(net364),
    .C(net347),
    .X(_1359_));
 sky130_fd_sc_hd__a221o_4 _3717_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ),
    .A2(net302),
    .B1(net345),
    .B2(net304),
    .C1(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__nand2_1 _3718_ (.A(_1358_),
    .B(_1360_),
    .Y(_1361_));
 sky130_fd_sc_hd__or2_1 _3719_ (.A(_1358_),
    .B(_1360_),
    .X(_1362_));
 sky130_fd_sc_hd__and2_1 _3720_ (.A(_1361_),
    .B(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__and2b_1 _3721_ (.A_N(net436),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[29] ),
    .X(_1364_));
 sky130_fd_sc_hd__a221o_1 _3722_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[29] ),
    .A2(net370),
    .B1(net367),
    .B2(net52),
    .C1(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__mux2_1 _3723_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[29] ),
    .A1(_1365_),
    .S(net372),
    .X(_1366_));
 sky130_fd_sc_hd__a22o_1 _3724_ (.A1(net2220),
    .A2(net307),
    .B1(net344),
    .B2(_1312_),
    .X(_1367_));
 sky130_fd_sc_hd__a21oi_4 _3725_ (.A1(net2198),
    .A2(net354),
    .B1(_1367_),
    .Y(_1368_));
 sky130_fd_sc_hd__nand2_1 _3726_ (.A(net377),
    .B(net2216),
    .Y(_1369_));
 sky130_fd_sc_hd__o21ai_4 _3727_ (.A1(net377),
    .A2(_1368_),
    .B1(_1369_),
    .Y(_1370_));
 sky130_fd_sc_hd__inv_2 _3728_ (.A(_1370_),
    .Y(_1371_));
 sky130_fd_sc_hd__and3_1 _3729_ (.A(net2198),
    .B(net365),
    .C(net348),
    .X(_1372_));
 sky130_fd_sc_hd__a221o_4 _3730_ (.A1(net2260),
    .A2(net303),
    .B1(net344),
    .B2(net305),
    .C1(_1372_),
    .X(_1373_));
 sky130_fd_sc_hd__or2_1 _3731_ (.A(_1370_),
    .B(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__nand2_1 _3732_ (.A(_1370_),
    .B(_1373_),
    .Y(_1375_));
 sky130_fd_sc_hd__and2_1 _3733_ (.A(_1374_),
    .B(_1375_),
    .X(_1376_));
 sky130_fd_sc_hd__a2111o_2 _3734_ (.A1(_1351_),
    .A2(_1352_),
    .B1(_1363_),
    .C1(_1376_),
    .D1(_1339_),
    .X(_1377_));
 sky130_fd_sc_hd__and2b_1 _3735_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[17] ),
    .X(_1378_));
 sky130_fd_sc_hd__a221o_2 _3736_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[17] ),
    .A2(net369),
    .B1(net366),
    .B2(net39),
    .C1(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__or2_2 _3737_ (.A(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[17] ),
    .B(net372),
    .X(_1380_));
 sky130_fd_sc_hd__o21ai_4 _3738_ (.A1(_1313_),
    .A2(_1379_),
    .B1(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__o21a_4 _3739_ (.A1(_1313_),
    .A2(_1379_),
    .B1(_1380_),
    .X(_1382_));
 sky130_fd_sc_hd__or3_1 _3740_ (.A(net354),
    .B(_1311_),
    .C(_1381_),
    .X(_1383_));
 sky130_fd_sc_hd__nand2_1 _3741_ (.A(net898),
    .B(net354),
    .Y(_1384_));
 sky130_fd_sc_hd__or3b_1 _3742_ (.A(net354),
    .B(net349),
    .C_N(net2253),
    .X(_1385_));
 sky130_fd_sc_hd__a31o_1 _3743_ (.A1(_1383_),
    .A2(_1384_),
    .A3(_1385_),
    .B1(net377),
    .X(_1386_));
 sky130_fd_sc_hd__nand2_1 _3744_ (.A(net377),
    .B(net2200),
    .Y(_1387_));
 sky130_fd_sc_hd__nand2_1 _3745_ (.A(_1386_),
    .B(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__and3_1 _3746_ (.A(net898),
    .B(net365),
    .C(net348),
    .X(_1389_));
 sky130_fd_sc_hd__a221oi_4 _3747_ (.A1(net2305),
    .A2(net303),
    .B1(_1382_),
    .B2(net305),
    .C1(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__a221o_2 _3748_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ),
    .A2(net303),
    .B1(_1382_),
    .B2(net305),
    .C1(_1389_),
    .X(_1391_));
 sky130_fd_sc_hd__nand3_1 _3749_ (.A(_1386_),
    .B(_1387_),
    .C(_1390_),
    .Y(_1392_));
 sky130_fd_sc_hd__a21o_1 _3750_ (.A1(_1386_),
    .A2(_1387_),
    .B1(_1390_),
    .X(_1393_));
 sky130_fd_sc_hd__and2b_1 _3751_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[19] ),
    .X(_1394_));
 sky130_fd_sc_hd__a221o_1 _3752_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[19] ),
    .A2(net369),
    .B1(net366),
    .B2(net41),
    .C1(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__mux2_1 _3753_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[19] ),
    .A1(_1395_),
    .S(net371),
    .X(_1396_));
 sky130_fd_sc_hd__and3_1 _3754_ (.A(net352),
    .B(net349),
    .C(net343),
    .X(_1397_));
 sky130_fd_sc_hd__a221o_1 _3755_ (.A1(net2168),
    .A2(net354),
    .B1(net307),
    .B2(net2204),
    .C1(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__mux2_2 _3756_ (.A0(net2132),
    .A1(_1398_),
    .S(net373),
    .X(_1399_));
 sky130_fd_sc_hd__and3_1 _3757_ (.A(net2168),
    .B(net364),
    .C(net347),
    .X(_1400_));
 sky130_fd_sc_hd__a221o_4 _3758_ (.A1(net2317),
    .A2(net302),
    .B1(net343),
    .B2(net304),
    .C1(_1400_),
    .X(_1401_));
 sky130_fd_sc_hd__or2_1 _3759_ (.A(_1399_),
    .B(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__nand2_1 _3760_ (.A(_1399_),
    .B(_1401_),
    .Y(_1403_));
 sky130_fd_sc_hd__and2_1 _3761_ (.A(_1402_),
    .B(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__and2b_1 _3762_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[16] ),
    .X(_1405_));
 sky130_fd_sc_hd__a221o_1 _3763_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[16] ),
    .A2(net369),
    .B1(net366),
    .B2(net38),
    .C1(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__mux2_1 _3764_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[16] ),
    .A1(_1406_),
    .S(net371),
    .X(_1407_));
 sky130_fd_sc_hd__and3_1 _3765_ (.A(net351),
    .B(net350),
    .C(net342),
    .X(_1408_));
 sky130_fd_sc_hd__a221oi_4 _3766_ (.A1(net2047),
    .A2(net353),
    .B1(net306),
    .B2(net2280),
    .C1(_1408_),
    .Y(_1409_));
 sky130_fd_sc_hd__inv_2 _3767_ (.A(_1409_),
    .Y(_1410_));
 sky130_fd_sc_hd__mux2_1 _3768_ (.A0(_1289_),
    .A1(_1409_),
    .S(net373),
    .X(_1411_));
 sky130_fd_sc_hd__mux2_1 _3769_ (.A0(net2075),
    .A1(_1410_),
    .S(net373),
    .X(_1412_));
 sky130_fd_sc_hd__and3_1 _3770_ (.A(net71),
    .B(net364),
    .C(net347),
    .X(_1413_));
 sky130_fd_sc_hd__a221o_4 _3771_ (.A1(net2303),
    .A2(net302),
    .B1(net342),
    .B2(net304),
    .C1(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__nand2_1 _3772_ (.A(_1412_),
    .B(_1414_),
    .Y(_1415_));
 sky130_fd_sc_hd__or2_1 _3773_ (.A(_1412_),
    .B(_1414_),
    .X(_1416_));
 sky130_fd_sc_hd__and2_1 _3774_ (.A(_1415_),
    .B(_1416_),
    .X(_1417_));
 sky130_fd_sc_hd__and2b_1 _3775_ (.A_N(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[18] ),
    .X(_1418_));
 sky130_fd_sc_hd__a221o_1 _3776_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[18] ),
    .A2(net370),
    .B1(net367),
    .B2(net40),
    .C1(_1418_),
    .X(_1419_));
 sky130_fd_sc_hd__mux2_1 _3777_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[18] ),
    .A1(_1419_),
    .S(net372),
    .X(_1420_));
 sky130_fd_sc_hd__and3_1 _3778_ (.A(net351),
    .B(net349),
    .C(net341),
    .X(_1421_));
 sky130_fd_sc_hd__a221o_2 _3779_ (.A1(net1977),
    .A2(net353),
    .B1(net306),
    .B2(net2292),
    .C1(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__mux2_4 _3780_ (.A0(net2148),
    .A1(_1422_),
    .S(net373),
    .X(_1423_));
 sky130_fd_sc_hd__and3_1 _3781_ (.A(net73),
    .B(net364),
    .C(net347),
    .X(_1424_));
 sky130_fd_sc_hd__a221o_4 _3782_ (.A1(net2347),
    .A2(net302),
    .B1(net341),
    .B2(net304),
    .C1(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__nand2_1 _3783_ (.A(_1423_),
    .B(_1425_),
    .Y(_1426_));
 sky130_fd_sc_hd__or2_1 _3784_ (.A(_1423_),
    .B(_1425_),
    .X(_1427_));
 sky130_fd_sc_hd__xor2_1 _3785_ (.A(_1423_),
    .B(_1425_),
    .X(_1428_));
 sky130_fd_sc_hd__a2111o_1 _3786_ (.A1(_1392_),
    .A2(_1393_),
    .B1(_1404_),
    .C1(_1417_),
    .D1(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__and2b_1 _3787_ (.A_N(net436),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[21] ),
    .X(_1430_));
 sky130_fd_sc_hd__a221o_1 _3788_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[21] ),
    .A2(net370),
    .B1(net367),
    .B2(net44),
    .C1(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__mux2_2 _3789_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[21] ),
    .A1(_1431_),
    .S(net372),
    .X(_1432_));
 sky130_fd_sc_hd__and3_1 _3790_ (.A(net352),
    .B(net349),
    .C(net340),
    .X(_1433_));
 sky130_fd_sc_hd__a221o_1 _3791_ (.A1(net2005),
    .A2(net354),
    .B1(net307),
    .B2(net2203),
    .C1(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__mux2_2 _3792_ (.A0(net2263),
    .A1(_1434_),
    .S(net374),
    .X(_1435_));
 sky130_fd_sc_hd__and3_1 _3793_ (.A(net2005),
    .B(net365),
    .C(net348),
    .X(_1436_));
 sky130_fd_sc_hd__a221o_4 _3794_ (.A1(net2310),
    .A2(net303),
    .B1(net340),
    .B2(net305),
    .C1(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__or2_1 _3795_ (.A(_1435_),
    .B(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__xor2_1 _3796_ (.A(_1435_),
    .B(_1437_),
    .X(_1439_));
 sky130_fd_sc_hd__and2b_1 _3797_ (.A_N(net436),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[22] ),
    .X(_1440_));
 sky130_fd_sc_hd__a221o_1 _3798_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[22] ),
    .A2(net370),
    .B1(net367),
    .B2(net45),
    .C1(_1440_),
    .X(_1441_));
 sky130_fd_sc_hd__mux2_4 _3799_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[22] ),
    .A1(_1441_),
    .S(net372),
    .X(_1442_));
 sky130_fd_sc_hd__and3_1 _3800_ (.A(net351),
    .B(net349),
    .C(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__a221o_4 _3801_ (.A1(net2185),
    .A2(net353),
    .B1(net306),
    .B2(net2316),
    .C1(_1443_),
    .X(_1444_));
 sky130_fd_sc_hd__mux2_2 _3802_ (.A0(net2181),
    .A1(_1444_),
    .S(net374),
    .X(_1445_));
 sky130_fd_sc_hd__and3_1 _3803_ (.A(net78),
    .B(net365),
    .C(net348),
    .X(_1446_));
 sky130_fd_sc_hd__a221o_4 _3804_ (.A1(net2293),
    .A2(net303),
    .B1(net339),
    .B2(net305),
    .C1(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__nand2_1 _3805_ (.A(_1445_),
    .B(net2294),
    .Y(_1448_));
 sky130_fd_sc_hd__xor2_1 _3806_ (.A(_1445_),
    .B(_1447_),
    .X(_1449_));
 sky130_fd_sc_hd__and2b_1 _3807_ (.A_N(net436),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[20] ),
    .X(_1450_));
 sky130_fd_sc_hd__a221o_1 _3808_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[20] ),
    .A2(net370),
    .B1(net367),
    .B2(net43),
    .C1(_1450_),
    .X(_1451_));
 sky130_fd_sc_hd__mux2_1 _3809_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[20] ),
    .A1(_1451_),
    .S(net372),
    .X(_1452_));
 sky130_fd_sc_hd__a22o_1 _3810_ (.A1(net2273),
    .A2(net307),
    .B1(net338),
    .B2(_1312_),
    .X(_1453_));
 sky130_fd_sc_hd__a21oi_4 _3811_ (.A1(net2080),
    .A2(net354),
    .B1(_1453_),
    .Y(_1454_));
 sky130_fd_sc_hd__nand2_1 _3812_ (.A(net377),
    .B(net2243),
    .Y(_1455_));
 sky130_fd_sc_hd__o21ai_4 _3813_ (.A1(net377),
    .A2(_1454_),
    .B1(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__and3_1 _3814_ (.A(net76),
    .B(net365),
    .C(net348),
    .X(_1457_));
 sky130_fd_sc_hd__a221o_4 _3815_ (.A1(net2333),
    .A2(net303),
    .B1(net338),
    .B2(net305),
    .C1(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__nand2_1 _3816_ (.A(_1456_),
    .B(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__or2_1 _3817_ (.A(_1456_),
    .B(_1458_),
    .X(_1460_));
 sky130_fd_sc_hd__and2b_1 _3818_ (.A_N(net436),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[23] ),
    .X(_1461_));
 sky130_fd_sc_hd__a221o_1 _3819_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[23] ),
    .A2(net370),
    .B1(net367),
    .B2(net46),
    .C1(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__mux2_1 _3820_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[23] ),
    .A1(_1462_),
    .S(net372),
    .X(_1463_));
 sky130_fd_sc_hd__and3_1 _3821_ (.A(net352),
    .B(net349),
    .C(net337),
    .X(_1464_));
 sky130_fd_sc_hd__a221o_1 _3822_ (.A1(net2016),
    .A2(net354),
    .B1(net307),
    .B2(net2266),
    .C1(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__mux2_2 _3823_ (.A0(net2210),
    .A1(_1465_),
    .S(net374),
    .X(_1466_));
 sky130_fd_sc_hd__and3_1 _3824_ (.A(net2016),
    .B(net365),
    .C(net348),
    .X(_1467_));
 sky130_fd_sc_hd__a221o_4 _3825_ (.A1(net2307),
    .A2(net303),
    .B1(net337),
    .B2(net305),
    .C1(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__or2_1 _3826_ (.A(_1466_),
    .B(_1468_),
    .X(_1469_));
 sky130_fd_sc_hd__xor2_1 _3827_ (.A(_1466_),
    .B(_1468_),
    .X(_1470_));
 sky130_fd_sc_hd__or3_1 _3828_ (.A(_1439_),
    .B(_1449_),
    .C(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__a21o_1 _3829_ (.A1(_1459_),
    .A2(_1460_),
    .B1(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__and2b_1 _3830_ (.A_N(net436),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[25] ),
    .X(_1473_));
 sky130_fd_sc_hd__a221o_1 _3831_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[25] ),
    .A2(net370),
    .B1(net367),
    .B2(net48),
    .C1(_1473_),
    .X(_1474_));
 sky130_fd_sc_hd__mux2_1 _3832_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[25] ),
    .A1(_1474_),
    .S(net372),
    .X(_1475_));
 sky130_fd_sc_hd__a22o_1 _3833_ (.A1(net2140),
    .A2(net307),
    .B1(net336),
    .B2(_1312_),
    .X(_1476_));
 sky130_fd_sc_hd__a21oi_4 _3834_ (.A1(net2006),
    .A2(net354),
    .B1(net2141),
    .Y(_1477_));
 sky130_fd_sc_hd__nand2_1 _3835_ (.A(net377),
    .B(net2281),
    .Y(_1478_));
 sky130_fd_sc_hd__o21ai_4 _3836_ (.A1(net377),
    .A2(_1477_),
    .B1(net2282),
    .Y(_1479_));
 sky130_fd_sc_hd__inv_2 _3837_ (.A(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__and3_1 _3838_ (.A(net2006),
    .B(net365),
    .C(net348),
    .X(_1481_));
 sky130_fd_sc_hd__a221o_4 _3839_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[25] ),
    .A2(net303),
    .B1(net336),
    .B2(net305),
    .C1(_1481_),
    .X(_1482_));
 sky130_fd_sc_hd__or2_1 _3840_ (.A(_1479_),
    .B(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__xor2_1 _3841_ (.A(_1479_),
    .B(_1482_),
    .X(_1484_));
 sky130_fd_sc_hd__and2b_1 _3842_ (.A_N(net436),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[26] ),
    .X(_1485_));
 sky130_fd_sc_hd__a221o_1 _3843_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[26] ),
    .A2(net370),
    .B1(net367),
    .B2(net49),
    .C1(_1485_),
    .X(_1486_));
 sky130_fd_sc_hd__mux2_2 _3844_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[26] ),
    .A1(_1486_),
    .S(net372),
    .X(_1487_));
 sky130_fd_sc_hd__and3_1 _3845_ (.A(net352),
    .B(net349),
    .C(net335),
    .X(_1488_));
 sky130_fd_sc_hd__a221o_2 _3846_ (.A1(net2143),
    .A2(net354),
    .B1(net307),
    .B2(net2208),
    .C1(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__mux2_2 _3847_ (.A0(net2233),
    .A1(_1489_),
    .S(net374),
    .X(_1490_));
 sky130_fd_sc_hd__and3_1 _3848_ (.A(net82),
    .B(net365),
    .C(net348),
    .X(_1491_));
 sky130_fd_sc_hd__a221o_4 _3849_ (.A1(net2342),
    .A2(net303),
    .B1(net335),
    .B2(net305),
    .C1(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__and2_1 _3850_ (.A(_1490_),
    .B(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__nor2_1 _3851_ (.A(_1490_),
    .B(_1492_),
    .Y(_1494_));
 sky130_fd_sc_hd__nor2_1 _3852_ (.A(_1493_),
    .B(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__and2b_1 _3853_ (.A_N(net436),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[24] ),
    .X(_1496_));
 sky130_fd_sc_hd__a221o_1 _3854_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[24] ),
    .A2(net370),
    .B1(net367),
    .B2(net47),
    .C1(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__mux2_8 _3855_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[24] ),
    .A1(_1497_),
    .S(net372),
    .X(_1498_));
 sky130_fd_sc_hd__a22o_1 _3856_ (.A1(net2291),
    .A2(net306),
    .B1(net334),
    .B2(_1312_),
    .X(_1499_));
 sky130_fd_sc_hd__a21oi_4 _3857_ (.A1(net2159),
    .A2(net355),
    .B1(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__nand2_1 _3858_ (.A(net377),
    .B(net2301),
    .Y(_1501_));
 sky130_fd_sc_hd__o21ai_4 _3859_ (.A1(net377),
    .A2(_1500_),
    .B1(_1501_),
    .Y(_1502_));
 sky130_fd_sc_hd__inv_2 _3860_ (.A(_1502_),
    .Y(_1503_));
 sky130_fd_sc_hd__and3_1 _3861_ (.A(net80),
    .B(net365),
    .C(net348),
    .X(_1504_));
 sky130_fd_sc_hd__a221o_4 _3862_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ),
    .A2(net303),
    .B1(net334),
    .B2(net305),
    .C1(_1504_),
    .X(_1505_));
 sky130_fd_sc_hd__nand2_1 _3863_ (.A(_1502_),
    .B(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hd__or2_1 _3864_ (.A(_1502_),
    .B(_1505_),
    .X(_1507_));
 sky130_fd_sc_hd__and2b_1 _3865_ (.A_N(net436),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[27] ),
    .X(_1508_));
 sky130_fd_sc_hd__a221o_1 _3866_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[27] ),
    .A2(net370),
    .B1(net367),
    .B2(net50),
    .C1(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__mux2_4 _3867_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[27] ),
    .A1(_1509_),
    .S(net372),
    .X(_1510_));
 sky130_fd_sc_hd__a22o_1 _3868_ (.A1(net2275),
    .A2(net306),
    .B1(net333),
    .B2(_1312_),
    .X(_1511_));
 sky130_fd_sc_hd__a21oi_4 _3869_ (.A1(net2178),
    .A2(net353),
    .B1(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__inv_2 _3870_ (.A(_1512_),
    .Y(_1513_));
 sky130_fd_sc_hd__mux2_4 _3871_ (.A0(net2186),
    .A1(_1513_),
    .S(net374),
    .X(_1514_));
 sky130_fd_sc_hd__and3_1 _3872_ (.A(net83),
    .B(net365),
    .C(net348),
    .X(_1515_));
 sky130_fd_sc_hd__a221o_4 _3873_ (.A1(net2330),
    .A2(net303),
    .B1(net333),
    .B2(net305),
    .C1(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__xor2_1 _3874_ (.A(_1514_),
    .B(_1516_),
    .X(_1517_));
 sky130_fd_sc_hd__a21o_1 _3875_ (.A1(_1506_),
    .A2(_1507_),
    .B1(_1484_),
    .X(_1518_));
 sky130_fd_sc_hd__or3_1 _3876_ (.A(_1495_),
    .B(_1517_),
    .C(_1518_),
    .X(_1519_));
 sky130_fd_sc_hd__or4_4 _3877_ (.A(_1377_),
    .B(_1429_),
    .C(_1472_),
    .D(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__and2b_1 _3878_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[3] ),
    .X(_1521_));
 sky130_fd_sc_hd__a221o_1 _3879_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[3] ),
    .A2(net369),
    .B1(net366),
    .B2(net56),
    .C1(_1521_),
    .X(_1522_));
 sky130_fd_sc_hd__mux2_2 _3880_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[3] ),
    .A1(_1522_),
    .S(net371),
    .X(_1523_));
 sky130_fd_sc_hd__and3_1 _3881_ (.A(net351),
    .B(net350),
    .C(net332),
    .X(_1524_));
 sky130_fd_sc_hd__a221oi_4 _3882_ (.A1(net1984),
    .A2(_1300_),
    .B1(net306),
    .B2(net2252),
    .C1(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__nand2_1 _3883_ (.A(net378),
    .B(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ),
    .Y(_1526_));
 sky130_fd_sc_hd__o21a_1 _3884_ (.A1(net378),
    .A2(_1525_),
    .B1(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__o21ai_2 _3885_ (.A1(net378),
    .A2(_1525_),
    .B1(_1526_),
    .Y(_1528_));
 sky130_fd_sc_hd__and3_1 _3886_ (.A(net89),
    .B(net364),
    .C(net347),
    .X(_1529_));
 sky130_fd_sc_hd__a221o_4 _3887_ (.A1(net2351),
    .A2(net302),
    .B1(net332),
    .B2(net304),
    .C1(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__or2_1 _3888_ (.A(net209),
    .B(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__xnor2_1 _3889_ (.A(net209),
    .B(_1530_),
    .Y(_1532_));
 sky130_fd_sc_hd__and2b_1 _3890_ (.A_N(net436),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[2] ),
    .X(_1533_));
 sky130_fd_sc_hd__a221o_1 _3891_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[2] ),
    .A2(net370),
    .B1(net367),
    .B2(net53),
    .C1(_1533_),
    .X(_1534_));
 sky130_fd_sc_hd__mux2_4 _3892_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[2] ),
    .A1(_1534_),
    .S(net372),
    .X(_1535_));
 sky130_fd_sc_hd__and3_1 _3893_ (.A(net352),
    .B(net349),
    .C(net331),
    .X(_1536_));
 sky130_fd_sc_hd__a221o_4 _3894_ (.A1(net860),
    .A2(net354),
    .B1(net307),
    .B2(net2325),
    .C1(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__and2_1 _3895_ (.A(net378),
    .B(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ),
    .X(_1538_));
 sky130_fd_sc_hd__a21oi_4 _3896_ (.A1(net373),
    .A2(_1537_),
    .B1(_1538_),
    .Y(_1539_));
 sky130_fd_sc_hd__a21o_1 _3897_ (.A1(net373),
    .A2(_1537_),
    .B1(_1538_),
    .X(_1540_));
 sky130_fd_sc_hd__and3_1 _3898_ (.A(net86),
    .B(net365),
    .C(net348),
    .X(_1541_));
 sky130_fd_sc_hd__a221o_4 _3899_ (.A1(net2298),
    .A2(net303),
    .B1(net331),
    .B2(net305),
    .C1(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__and2_1 _3900_ (.A(net203),
    .B(_1542_),
    .X(_1543_));
 sky130_fd_sc_hd__nor2_1 _3901_ (.A(net203),
    .B(_1542_),
    .Y(_1544_));
 sky130_fd_sc_hd__xnor2_1 _3902_ (.A(net203),
    .B(_1542_),
    .Y(_1545_));
 sky130_fd_sc_hd__nand2_1 _3903_ (.A(_1532_),
    .B(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hd__a22o_1 _3904_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[1] ),
    .A2(net369),
    .B1(net366),
    .B2(net42),
    .X(_1547_));
 sky130_fd_sc_hd__a21o_4 _3905_ (.A1(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[1] ),
    .A2(_1313_),
    .B1(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__and3_1 _3906_ (.A(net352),
    .B(net349),
    .C(net330),
    .X(_1549_));
 sky130_fd_sc_hd__nor2_1 _3907_ (.A(_1290_),
    .B(net352),
    .Y(_1550_));
 sky130_fd_sc_hd__and3_2 _3908_ (.A(net2335),
    .B(net351),
    .C(_1311_),
    .X(_1551_));
 sky130_fd_sc_hd__o31a_1 _3909_ (.A1(_1549_),
    .A2(_1550_),
    .A3(_1551_),
    .B1(net373),
    .X(_1552_));
 sky130_fd_sc_hd__nand2_1 _3910_ (.A(net378),
    .B(net2136),
    .Y(_1553_));
 sky130_fd_sc_hd__inv_2 _3911_ (.A(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__nor2_2 _3912_ (.A(_1552_),
    .B(_1554_),
    .Y(_1555_));
 sky130_fd_sc_hd__or2_1 _3913_ (.A(_1552_),
    .B(_1554_),
    .X(_1556_));
 sky130_fd_sc_hd__and3_1 _3914_ (.A(net2066),
    .B(net364),
    .C(net347),
    .X(_1557_));
 sky130_fd_sc_hd__a221o_4 _3915_ (.A1(net2350),
    .A2(net302),
    .B1(net330),
    .B2(net304),
    .C1(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__inv_2 _3916_ (.A(_1558_),
    .Y(_1559_));
 sky130_fd_sc_hd__or2_1 _3917_ (.A(net198),
    .B(_1558_),
    .X(_1560_));
 sky130_fd_sc_hd__nand2_1 _3918_ (.A(net198),
    .B(_1558_),
    .Y(_1561_));
 sky130_fd_sc_hd__and2_1 _3919_ (.A(_1560_),
    .B(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__a22o_1 _3920_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[0] ),
    .A2(net369),
    .B1(net366),
    .B2(net31),
    .X(_1563_));
 sky130_fd_sc_hd__a21o_2 _3921_ (.A1(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[0] ),
    .A2(_1313_),
    .B1(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__and3_1 _3922_ (.A(net351),
    .B(net349),
    .C(net329),
    .X(_1565_));
 sky130_fd_sc_hd__a221o_2 _3923_ (.A1(net2007),
    .A2(net353),
    .B1(net306),
    .B2(net2236),
    .C1(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__mux2_1 _3924_ (.A0(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[0] ),
    .A1(_1566_),
    .S(net373),
    .X(_1567_));
 sky130_fd_sc_hd__and3_1 _3925_ (.A(net64),
    .B(net364),
    .C(net347),
    .X(_1568_));
 sky130_fd_sc_hd__a221o_4 _3926_ (.A1(net2300),
    .A2(net302),
    .B1(net329),
    .B2(net304),
    .C1(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__inv_2 _3927_ (.A(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__nand2_2 _3928_ (.A(net194),
    .B(_1569_),
    .Y(_1571_));
 sky130_fd_sc_hd__or2_1 _3929_ (.A(net194),
    .B(_1569_),
    .X(_1572_));
 sky130_fd_sc_hd__and2b_1 _3930_ (.A_N(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[7] ),
    .X(_1573_));
 sky130_fd_sc_hd__a221o_2 _3931_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[7] ),
    .A2(net369),
    .B1(net366),
    .B2(net60),
    .C1(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__mux2_1 _3932_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[7] ),
    .A1(_1574_),
    .S(net371),
    .X(_1575_));
 sky130_fd_sc_hd__and3_1 _3933_ (.A(net351),
    .B(net349),
    .C(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__a221o_2 _3934_ (.A1(net2034),
    .A2(net353),
    .B1(net307),
    .B2(net2250),
    .C1(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__mux2_4 _3935_ (.A0(net2160),
    .A1(_1577_),
    .S(net373),
    .X(_1578_));
 sky130_fd_sc_hd__and3_1 _3936_ (.A(net93),
    .B(net364),
    .C(net347),
    .X(_1579_));
 sky130_fd_sc_hd__a221o_4 _3937_ (.A1(net2320),
    .A2(net302),
    .B1(net328),
    .B2(net304),
    .C1(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__xor2_1 _3938_ (.A(_1578_),
    .B(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__and2b_1 _3939_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[4] ),
    .X(_1582_));
 sky130_fd_sc_hd__a221o_1 _3940_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[4] ),
    .A2(net369),
    .B1(net366),
    .B2(net57),
    .C1(_1582_),
    .X(_1583_));
 sky130_fd_sc_hd__mux2_2 _3941_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[4] ),
    .A1(_1583_),
    .S(net371),
    .X(_1584_));
 sky130_fd_sc_hd__and3_1 _3942_ (.A(net351),
    .B(net350),
    .C(net327),
    .X(_1585_));
 sky130_fd_sc_hd__a221o_4 _3943_ (.A1(net1928),
    .A2(net353),
    .B1(net306),
    .B2(net2299),
    .C1(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__and2_1 _3944_ (.A(net378),
    .B(net2229),
    .X(_1587_));
 sky130_fd_sc_hd__a21oi_1 _3945_ (.A1(net373),
    .A2(_1586_),
    .B1(_1587_),
    .Y(_1588_));
 sky130_fd_sc_hd__a21o_2 _3946_ (.A1(net373),
    .A2(_1586_),
    .B1(_1587_),
    .X(_1589_));
 sky130_fd_sc_hd__and3_1 _3947_ (.A(net1928),
    .B(net365),
    .C(net348),
    .X(_1590_));
 sky130_fd_sc_hd__a221o_4 _3948_ (.A1(net2349),
    .A2(net302),
    .B1(net327),
    .B2(net304),
    .C1(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__nand2_1 _3949_ (.A(net187),
    .B(_1591_),
    .Y(_1592_));
 sky130_fd_sc_hd__or2_1 _3950_ (.A(net187),
    .B(_1591_),
    .X(_1593_));
 sky130_fd_sc_hd__and2b_1 _3951_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[6] ),
    .X(_1594_));
 sky130_fd_sc_hd__a221o_1 _3952_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[6] ),
    .A2(net369),
    .B1(net366),
    .B2(net59),
    .C1(_1594_),
    .X(_1595_));
 sky130_fd_sc_hd__mux2_2 _3953_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[6] ),
    .A1(_1595_),
    .S(net371),
    .X(_1596_));
 sky130_fd_sc_hd__and3_1 _3954_ (.A(net352),
    .B(net349),
    .C(net326),
    .X(_1597_));
 sky130_fd_sc_hd__a221o_4 _3955_ (.A1(net2067),
    .A2(_1300_),
    .B1(net307),
    .B2(net2268),
    .C1(_1597_),
    .X(_1598_));
 sky130_fd_sc_hd__mux2_4 _3956_ (.A0(net2175),
    .A1(_1598_),
    .S(net373),
    .X(_1599_));
 sky130_fd_sc_hd__and3_1 _3957_ (.A(net92),
    .B(net364),
    .C(net347),
    .X(_1600_));
 sky130_fd_sc_hd__a221o_4 _3958_ (.A1(net2329),
    .A2(net303),
    .B1(net326),
    .B2(net305),
    .C1(_1600_),
    .X(_1601_));
 sky130_fd_sc_hd__nand2_1 _3959_ (.A(_1599_),
    .B(_1601_),
    .Y(_1602_));
 sky130_fd_sc_hd__xor2_1 _3960_ (.A(_1599_),
    .B(_1601_),
    .X(_1603_));
 sky130_fd_sc_hd__and2b_1 _3961_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[5] ),
    .X(_1604_));
 sky130_fd_sc_hd__a221o_2 _3962_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[5] ),
    .A2(net370),
    .B1(net367),
    .B2(net58),
    .C1(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__or2_2 _3963_ (.A(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[5] ),
    .B(net371),
    .X(_1606_));
 sky130_fd_sc_hd__o21ai_4 _3964_ (.A1(_1313_),
    .A2(_1605_),
    .B1(_1606_),
    .Y(_1607_));
 sky130_fd_sc_hd__o21a_4 _3965_ (.A1(_1313_),
    .A2(_1605_),
    .B1(_1606_),
    .X(_1608_));
 sky130_fd_sc_hd__and3_1 _3966_ (.A(net351),
    .B(net350),
    .C(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__and2_1 _3967_ (.A(net2152),
    .B(net353),
    .X(_1610_));
 sky130_fd_sc_hd__and3_1 _3968_ (.A(net2209),
    .B(net351),
    .C(_1311_),
    .X(_1611_));
 sky130_fd_sc_hd__o31a_2 _3969_ (.A1(_1609_),
    .A2(_1610_),
    .A3(_1611_),
    .B1(net374),
    .X(_1612_));
 sky130_fd_sc_hd__and2_1 _3970_ (.A(net378),
    .B(net2170),
    .X(_1613_));
 sky130_fd_sc_hd__or2_1 _3971_ (.A(_1612_),
    .B(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__and3_1 _3972_ (.A(net91),
    .B(net365),
    .C(net348),
    .X(_1615_));
 sky130_fd_sc_hd__a221o_4 _3973_ (.A1(net2340),
    .A2(net302),
    .B1(_1608_),
    .B2(net304),
    .C1(_1615_),
    .X(_1616_));
 sky130_fd_sc_hd__or3_1 _3974_ (.A(_1612_),
    .B(_1613_),
    .C(_1616_),
    .X(_1617_));
 sky130_fd_sc_hd__o21ai_1 _3975_ (.A1(_1612_),
    .A2(_1613_),
    .B1(_1616_),
    .Y(_1618_));
 sky130_fd_sc_hd__and2_1 _3976_ (.A(_1617_),
    .B(_1618_),
    .X(_1619_));
 sky130_fd_sc_hd__a2111o_1 _3977_ (.A1(_1592_),
    .A2(_1593_),
    .B1(_1603_),
    .C1(_1619_),
    .D1(_1581_),
    .X(_1620_));
 sky130_fd_sc_hd__a2111o_1 _3978_ (.A1(_1571_),
    .A2(_1572_),
    .B1(_1620_),
    .C1(_1562_),
    .D1(_1546_),
    .X(_1621_));
 sky130_fd_sc_hd__and2b_1 _3979_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[9] ),
    .X(_1622_));
 sky130_fd_sc_hd__a221o_1 _3980_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[9] ),
    .A2(net369),
    .B1(net366),
    .B2(net62),
    .C1(_1622_),
    .X(_1623_));
 sky130_fd_sc_hd__mux2_2 _3981_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[9] ),
    .A1(_1623_),
    .S(net371),
    .X(_1624_));
 sky130_fd_sc_hd__and3_1 _3982_ (.A(net351),
    .B(net350),
    .C(net325),
    .X(_1625_));
 sky130_fd_sc_hd__a221o_2 _3983_ (.A1(net2104),
    .A2(net353),
    .B1(net306),
    .B2(net2344),
    .C1(_1625_),
    .X(_1626_));
 sky130_fd_sc_hd__mux2_4 _3984_ (.A0(net2240),
    .A1(_1626_),
    .S(net373),
    .X(_1627_));
 sky130_fd_sc_hd__and3_1 _3985_ (.A(net95),
    .B(net364),
    .C(net347),
    .X(_1628_));
 sky130_fd_sc_hd__a221o_4 _3986_ (.A1(net2336),
    .A2(net302),
    .B1(net325),
    .B2(net304),
    .C1(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__xor2_1 _3987_ (.A(_1627_),
    .B(_1629_),
    .X(_1630_));
 sky130_fd_sc_hd__and2b_1 _3988_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[10] ),
    .X(_1631_));
 sky130_fd_sc_hd__a221o_1 _3989_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[10] ),
    .A2(net369),
    .B1(net366),
    .B2(net32),
    .C1(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__mux2_2 _3990_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[10] ),
    .A1(_1632_),
    .S(net371),
    .X(_1633_));
 sky130_fd_sc_hd__and3_1 _3991_ (.A(net351),
    .B(net350),
    .C(net324),
    .X(_1634_));
 sky130_fd_sc_hd__a221o_4 _3992_ (.A1(net962),
    .A2(net353),
    .B1(net306),
    .B2(net2223),
    .C1(_1634_),
    .X(_1635_));
 sky130_fd_sc_hd__mux2_4 _3993_ (.A0(net2189),
    .A1(_1635_),
    .S(net374),
    .X(_1636_));
 sky130_fd_sc_hd__and3_1 _3994_ (.A(net65),
    .B(_1323_),
    .C(_1327_),
    .X(_1637_));
 sky130_fd_sc_hd__a221o_4 _3995_ (.A1(net2346),
    .A2(_1336_),
    .B1(net324),
    .B2(_1334_),
    .C1(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__nand2_1 _3996_ (.A(_1636_),
    .B(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__or2_1 _3997_ (.A(_1636_),
    .B(_1638_),
    .X(_1640_));
 sky130_fd_sc_hd__xor2_1 _3998_ (.A(_1636_),
    .B(_1638_),
    .X(_1641_));
 sky130_fd_sc_hd__and2b_1 _3999_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[8] ),
    .X(_1642_));
 sky130_fd_sc_hd__a221o_1 _4000_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[8] ),
    .A2(net370),
    .B1(net367),
    .B2(net61),
    .C1(_1642_),
    .X(_1643_));
 sky130_fd_sc_hd__mux2_1 _4001_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[8] ),
    .A1(_1643_),
    .S(net371),
    .X(_1644_));
 sky130_fd_sc_hd__a22o_1 _4002_ (.A1(net2256),
    .A2(net306),
    .B1(net323),
    .B2(_1312_),
    .X(_1645_));
 sky130_fd_sc_hd__a21oi_4 _4003_ (.A1(net2008),
    .A2(net353),
    .B1(net2257),
    .Y(_1646_));
 sky130_fd_sc_hd__nand2_1 _4004_ (.A(net377),
    .B(net2224),
    .Y(_1647_));
 sky130_fd_sc_hd__o21ai_4 _4005_ (.A1(net377),
    .A2(_1646_),
    .B1(_1647_),
    .Y(_1648_));
 sky130_fd_sc_hd__and3_1 _4006_ (.A(net94),
    .B(_1323_),
    .C(_1327_),
    .X(_1649_));
 sky130_fd_sc_hd__a221o_4 _4007_ (.A1(net2339),
    .A2(net302),
    .B1(net323),
    .B2(net304),
    .C1(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__nand2_1 _4008_ (.A(_1648_),
    .B(_1650_),
    .Y(_1651_));
 sky130_fd_sc_hd__or2_1 _4009_ (.A(_1648_),
    .B(_1650_),
    .X(_1652_));
 sky130_fd_sc_hd__and2b_1 _4010_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[11] ),
    .X(_1653_));
 sky130_fd_sc_hd__a221o_1 _4011_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[11] ),
    .A2(net369),
    .B1(net366),
    .B2(net33),
    .C1(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__mux2_2 _4012_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[11] ),
    .A1(_1654_),
    .S(net371),
    .X(_1655_));
 sky130_fd_sc_hd__and3_1 _4013_ (.A(net352),
    .B(net349),
    .C(net322),
    .X(_1656_));
 sky130_fd_sc_hd__a221o_2 _4014_ (.A1(net778),
    .A2(net354),
    .B1(net307),
    .B2(net2276),
    .C1(_1656_),
    .X(_1657_));
 sky130_fd_sc_hd__mux2_4 _4015_ (.A0(net2214),
    .A1(_1657_),
    .S(net374),
    .X(_1658_));
 sky130_fd_sc_hd__and3_1 _4016_ (.A(net66),
    .B(net364),
    .C(net347),
    .X(_1659_));
 sky130_fd_sc_hd__a221o_4 _4017_ (.A1(net2341),
    .A2(net302),
    .B1(net322),
    .B2(net304),
    .C1(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__or2_1 _4018_ (.A(_1658_),
    .B(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__xor2_1 _4019_ (.A(_1658_),
    .B(_1660_),
    .X(_1662_));
 sky130_fd_sc_hd__or3_1 _4020_ (.A(_1630_),
    .B(_1641_),
    .C(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__a21o_1 _4021_ (.A1(_1651_),
    .A2(_1652_),
    .B1(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__and2b_1 _4022_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[13] ),
    .X(_1665_));
 sky130_fd_sc_hd__a221o_1 _4023_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[13] ),
    .A2(net369),
    .B1(net366),
    .B2(net35),
    .C1(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__mux2_1 _4024_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[13] ),
    .A1(_1666_),
    .S(net371),
    .X(_1667_));
 sky130_fd_sc_hd__and3_1 _4025_ (.A(net351),
    .B(net349),
    .C(net321),
    .X(_1668_));
 sky130_fd_sc_hd__a221o_4 _4026_ (.A1(net1855),
    .A2(net353),
    .B1(net306),
    .B2(net2269),
    .C1(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__mux2_2 _4027_ (.A0(net2199),
    .A1(_1669_),
    .S(net373),
    .X(_1670_));
 sky130_fd_sc_hd__inv_2 _4028_ (.A(_1670_),
    .Y(_1671_));
 sky130_fd_sc_hd__and3_1 _4029_ (.A(net68),
    .B(net364),
    .C(net347),
    .X(_1672_));
 sky130_fd_sc_hd__a221o_4 _4030_ (.A1(net2314),
    .A2(net302),
    .B1(net321),
    .B2(net304),
    .C1(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__or2_1 _4031_ (.A(_1670_),
    .B(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__nand2_1 _4032_ (.A(_1670_),
    .B(_1673_),
    .Y(_1675_));
 sky130_fd_sc_hd__and2_1 _4033_ (.A(_1674_),
    .B(_1675_),
    .X(_1676_));
 sky130_fd_sc_hd__and2b_1 _4034_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[14] ),
    .X(_1677_));
 sky130_fd_sc_hd__a221o_1 _4035_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[14] ),
    .A2(net369),
    .B1(net366),
    .B2(net36),
    .C1(_1677_),
    .X(_1678_));
 sky130_fd_sc_hd__mux2_1 _4036_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[14] ),
    .A1(_1678_),
    .S(net371),
    .X(_1679_));
 sky130_fd_sc_hd__and3_1 _4037_ (.A(net351),
    .B(net350),
    .C(net320),
    .X(_1680_));
 sky130_fd_sc_hd__a221o_4 _4038_ (.A1(net2147),
    .A2(net353),
    .B1(net306),
    .B2(net2255),
    .C1(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__mux2_2 _4039_ (.A0(net2193),
    .A1(_1681_),
    .S(net373),
    .X(_1682_));
 sky130_fd_sc_hd__and3_1 _4040_ (.A(net2147),
    .B(net364),
    .C(net347),
    .X(_1683_));
 sky130_fd_sc_hd__a221o_4 _4041_ (.A1(net2321),
    .A2(_1336_),
    .B1(net320),
    .B2(_1334_),
    .C1(_1683_),
    .X(_1684_));
 sky130_fd_sc_hd__nand2_1 _4042_ (.A(_1682_),
    .B(_1684_),
    .Y(_1685_));
 sky130_fd_sc_hd__or2_1 _4043_ (.A(_1682_),
    .B(_1684_),
    .X(_1686_));
 sky130_fd_sc_hd__and2_1 _4044_ (.A(_1685_),
    .B(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__and2b_1 _4045_ (.A_N(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[12] ),
    .X(_1688_));
 sky130_fd_sc_hd__a221o_1 _4046_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[12] ),
    .A2(net370),
    .B1(net367),
    .B2(net34),
    .C1(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__mux2_2 _4047_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[12] ),
    .A1(_1689_),
    .S(net371),
    .X(_1690_));
 sky130_fd_sc_hd__a22o_1 _4048_ (.A1(net2145),
    .A2(net306),
    .B1(net319),
    .B2(_1312_),
    .X(_1691_));
 sky130_fd_sc_hd__a21oi_4 _4049_ (.A1(net2130),
    .A2(net353),
    .B1(net2146),
    .Y(_1692_));
 sky130_fd_sc_hd__nand2_1 _4050_ (.A(net378),
    .B(net2164),
    .Y(_1693_));
 sky130_fd_sc_hd__o21ai_4 _4051_ (.A1(net378),
    .A2(_1692_),
    .B1(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__inv_2 _4052_ (.A(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__and3_1 _4053_ (.A(net67),
    .B(net364),
    .C(net347),
    .X(_1696_));
 sky130_fd_sc_hd__a221o_4 _4054_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ),
    .A2(net302),
    .B1(net319),
    .B2(net304),
    .C1(_1696_),
    .X(_1697_));
 sky130_fd_sc_hd__nand2_1 _4055_ (.A(_1694_),
    .B(_1697_),
    .Y(_1698_));
 sky130_fd_sc_hd__or2_1 _4056_ (.A(_1694_),
    .B(_1697_),
    .X(_1699_));
 sky130_fd_sc_hd__and2b_1 _4057_ (.A_N(net435),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[15] ),
    .X(_1700_));
 sky130_fd_sc_hd__a221o_1 _4058_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[15] ),
    .A2(net369),
    .B1(net366),
    .B2(net37),
    .C1(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__mux2_2 _4059_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[15] ),
    .A1(_1701_),
    .S(net371),
    .X(_1702_));
 sky130_fd_sc_hd__and3_1 _4060_ (.A(net351),
    .B(net350),
    .C(net318),
    .X(_1703_));
 sky130_fd_sc_hd__a221o_4 _4061_ (.A1(net2129),
    .A2(net353),
    .B1(net306),
    .B2(net2279),
    .C1(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__mux2_2 _4062_ (.A0(net2226),
    .A1(_1704_),
    .S(net373),
    .X(_1705_));
 sky130_fd_sc_hd__and3_1 _4063_ (.A(net70),
    .B(_1323_),
    .C(_1327_),
    .X(_1706_));
 sky130_fd_sc_hd__a221o_4 _4064_ (.A1(net2343),
    .A2(net302),
    .B1(net318),
    .B2(net304),
    .C1(_1706_),
    .X(_1707_));
 sky130_fd_sc_hd__or2_1 _4065_ (.A(_1705_),
    .B(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__nand2_1 _4066_ (.A(_1705_),
    .B(_1707_),
    .Y(_1709_));
 sky130_fd_sc_hd__and2_1 _4067_ (.A(_1708_),
    .B(_1709_),
    .X(_1710_));
 sky130_fd_sc_hd__or3_1 _4068_ (.A(_1676_),
    .B(_1687_),
    .C(_1710_),
    .X(_1711_));
 sky130_fd_sc_hd__a21o_1 _4069_ (.A1(_1698_),
    .A2(_1699_),
    .B1(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__or4_4 _4070_ (.A(_1520_),
    .B(_1621_),
    .C(_1664_),
    .D(_1712_),
    .X(_1713_));
 sky130_fd_sc_hd__nand2b_1 _4071_ (.A_N(_1601_),
    .B(_1599_),
    .Y(_1714_));
 sky130_fd_sc_hd__nand2b_1 _4072_ (.A_N(_1616_),
    .B(_1614_),
    .Y(_1715_));
 sky130_fd_sc_hd__a211o_1 _4073_ (.A1(_1617_),
    .A2(_1618_),
    .B1(net190),
    .C1(_1591_),
    .X(_1716_));
 sky130_fd_sc_hd__a21o_1 _4074_ (.A1(_1715_),
    .A2(_1716_),
    .B1(_1603_),
    .X(_1717_));
 sky130_fd_sc_hd__a21o_1 _4075_ (.A1(_1714_),
    .A2(_1717_),
    .B1(_1581_),
    .X(_1718_));
 sky130_fd_sc_hd__nand2b_1 _4076_ (.A_N(_1580_),
    .B(_1578_),
    .Y(_1719_));
 sky130_fd_sc_hd__o21a_1 _4077_ (.A1(net195),
    .A2(_1570_),
    .B1(net198),
    .X(_1720_));
 sky130_fd_sc_hd__or3_2 _4078_ (.A(net198),
    .B(net195),
    .C(_1570_),
    .X(_1721_));
 sky130_fd_sc_hd__inv_2 _4079_ (.A(_1721_),
    .Y(_1722_));
 sky130_fd_sc_hd__o2111ai_1 _4080_ (.A1(_1559_),
    .A2(_1720_),
    .B1(_1721_),
    .C1(_1545_),
    .D1(_1532_),
    .Y(_1723_));
 sky130_fd_sc_hd__or2_1 _4081_ (.A(net214),
    .B(_1530_),
    .X(_1724_));
 sky130_fd_sc_hd__or3b_1 _4082_ (.A(_1542_),
    .B(net206),
    .C_N(_1532_),
    .X(_1725_));
 sky130_fd_sc_hd__a31o_1 _4083_ (.A1(_1723_),
    .A2(_1724_),
    .A3(_1725_),
    .B1(_1620_),
    .X(_1726_));
 sky130_fd_sc_hd__a31o_1 _4084_ (.A1(_1718_),
    .A2(_1719_),
    .A3(_1726_),
    .B1(_1664_),
    .X(_1727_));
 sky130_fd_sc_hd__nand2b_1 _4085_ (.A_N(_1638_),
    .B(_1636_),
    .Y(_1728_));
 sky130_fd_sc_hd__nand2b_1 _4086_ (.A_N(_1629_),
    .B(_1627_),
    .Y(_1729_));
 sky130_fd_sc_hd__or3b_1 _4087_ (.A(_1630_),
    .B(_1650_),
    .C_N(_1648_),
    .X(_1730_));
 sky130_fd_sc_hd__a21o_1 _4088_ (.A1(_1729_),
    .A2(_1730_),
    .B1(_1641_),
    .X(_1731_));
 sky130_fd_sc_hd__a21o_1 _4089_ (.A1(_1728_),
    .A2(_1731_),
    .B1(_1662_),
    .X(_1732_));
 sky130_fd_sc_hd__nand2b_1 _4090_ (.A_N(_1660_),
    .B(_1658_),
    .Y(_1733_));
 sky130_fd_sc_hd__a31o_1 _4091_ (.A1(_1727_),
    .A2(_1732_),
    .A3(_1733_),
    .B1(_1712_),
    .X(_1734_));
 sky130_fd_sc_hd__nand2b_1 _4092_ (.A_N(_1684_),
    .B(_1682_),
    .Y(_1735_));
 sky130_fd_sc_hd__o32a_1 _4093_ (.A1(_1676_),
    .A2(_1695_),
    .A3(_1697_),
    .B1(_1673_),
    .B2(_1671_),
    .X(_1736_));
 sky130_fd_sc_hd__o21a_1 _4094_ (.A1(_1687_),
    .A2(_1736_),
    .B1(_1735_),
    .X(_1737_));
 sky130_fd_sc_hd__or2_1 _4095_ (.A(_1710_),
    .B(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__nand2b_1 _4096_ (.A_N(_1707_),
    .B(_1705_),
    .Y(_1739_));
 sky130_fd_sc_hd__a31oi_1 _4097_ (.A1(_1734_),
    .A2(_1738_),
    .A3(_1739_),
    .B1(_1520_),
    .Y(_1740_));
 sky130_fd_sc_hd__nand2_1 _4098_ (.A(_1321_),
    .B(_1338_),
    .Y(_1741_));
 sky130_fd_sc_hd__nand2b_1 _4099_ (.A_N(_1360_),
    .B(_1358_),
    .Y(_1742_));
 sky130_fd_sc_hd__o32a_1 _4100_ (.A1(_1348_),
    .A2(_1350_),
    .A3(_1376_),
    .B1(_1373_),
    .B2(_1371_),
    .X(_1743_));
 sky130_fd_sc_hd__o21a_1 _4101_ (.A1(_1363_),
    .A2(_1743_),
    .B1(_1742_),
    .X(_1744_));
 sky130_fd_sc_hd__o21ai_4 _4102_ (.A1(_1339_),
    .A2(_1744_),
    .B1(_1741_),
    .Y(_1745_));
 sky130_fd_sc_hd__nand2b_1 _4103_ (.A_N(_1401_),
    .B(_1399_),
    .Y(_1746_));
 sky130_fd_sc_hd__nand2b_1 _4104_ (.A_N(_1425_),
    .B(_1423_),
    .Y(_1747_));
 sky130_fd_sc_hd__and2_1 _4105_ (.A(_1388_),
    .B(_1390_),
    .X(_1748_));
 sky130_fd_sc_hd__a211oi_1 _4106_ (.A1(_1392_),
    .A2(_1393_),
    .B1(_1411_),
    .C1(_1414_),
    .Y(_1749_));
 sky130_fd_sc_hd__o21bai_1 _4107_ (.A1(_1748_),
    .A2(_1749_),
    .B1_N(_1428_),
    .Y(_1750_));
 sky130_fd_sc_hd__a21o_1 _4108_ (.A1(_1747_),
    .A2(_1750_),
    .B1(_1404_),
    .X(_1751_));
 sky130_fd_sc_hd__a21o_1 _4109_ (.A1(_1746_),
    .A2(_1751_),
    .B1(_1472_),
    .X(_1752_));
 sky130_fd_sc_hd__nand2b_1 _4110_ (.A_N(_1447_),
    .B(_1445_),
    .Y(_1753_));
 sky130_fd_sc_hd__nand2b_1 _4111_ (.A_N(_1437_),
    .B(_1435_),
    .Y(_1754_));
 sky130_fd_sc_hd__or3b_1 _4112_ (.A(_1439_),
    .B(_1458_),
    .C_N(_1456_),
    .X(_1755_));
 sky130_fd_sc_hd__a21o_1 _4113_ (.A1(_1754_),
    .A2(_1755_),
    .B1(_1449_),
    .X(_1756_));
 sky130_fd_sc_hd__a21o_1 _4114_ (.A1(_1753_),
    .A2(_1756_),
    .B1(_1470_),
    .X(_1757_));
 sky130_fd_sc_hd__nand2b_1 _4115_ (.A_N(_1468_),
    .B(_1466_),
    .Y(_1758_));
 sky130_fd_sc_hd__a31o_1 _4116_ (.A1(_1752_),
    .A2(_1757_),
    .A3(_1758_),
    .B1(_1519_),
    .X(_1759_));
 sky130_fd_sc_hd__nand2b_1 _4117_ (.A_N(_1492_),
    .B(_1490_),
    .Y(_1760_));
 sky130_fd_sc_hd__o32a_1 _4118_ (.A1(_1484_),
    .A2(_1503_),
    .A3(_1505_),
    .B1(_1482_),
    .B2(_1480_),
    .X(_1761_));
 sky130_fd_sc_hd__o21a_1 _4119_ (.A1(_1495_),
    .A2(_1761_),
    .B1(_1760_),
    .X(_1762_));
 sky130_fd_sc_hd__or2_1 _4120_ (.A(_1517_),
    .B(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__nand2b_1 _4121_ (.A_N(_1516_),
    .B(_1514_),
    .Y(_1764_));
 sky130_fd_sc_hd__a31oi_4 _4122_ (.A1(_1759_),
    .A2(_1763_),
    .A3(_1764_),
    .B1(_1377_),
    .Y(_1765_));
 sky130_fd_sc_hd__o31ai_2 _4123_ (.A1(_1740_),
    .A2(_1745_),
    .A3(_1765_),
    .B1(_1713_),
    .Y(_1766_));
 sky130_fd_sc_hd__nand2_1 _4124_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ),
    .Y(_1767_));
 sky130_fd_sc_hd__xor2_1 _4125_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .B(_1766_),
    .X(_1768_));
 sky130_fd_sc_hd__and3b_2 _4126_ (.A_N(net2231),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .C(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .X(_1769_));
 sky130_fd_sc_hd__inv_2 _4127_ (.A(_1769_),
    .Y(_1770_));
 sky130_fd_sc_hd__nand2b_4 _4128_ (.A_N(net2354),
    .B(net2323),
    .Y(_1771_));
 sky130_fd_sc_hd__nand2b_4 _4129_ (.A_N(net2323),
    .B(net2326),
    .Y(_1772_));
 sky130_fd_sc_hd__or3_4 _4130_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .C(net2231),
    .X(_1773_));
 sky130_fd_sc_hd__o22a_1 _4131_ (.A1(_1770_),
    .A2(net2324),
    .B1(_1772_),
    .B2(_1773_),
    .X(_1774_));
 sky130_fd_sc_hd__or3b_4 _4132_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .B(net2287),
    .C_N(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .X(_1775_));
 sky130_fd_sc_hd__o21a_1 _4133_ (.A1(_1772_),
    .A2(_1775_),
    .B1(_1774_),
    .X(_1776_));
 sky130_fd_sc_hd__or2_1 _4134_ (.A(_1770_),
    .B(_1772_),
    .X(_1777_));
 sky130_fd_sc_hd__mux2_1 _4135_ (.A0(_1776_),
    .A1(_1777_),
    .S(_1713_),
    .X(_1778_));
 sky130_fd_sc_hd__o31ai_1 _4136_ (.A1(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .A2(_1767_),
    .A3(_1768_),
    .B1(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hd__a21oi_1 _4137_ (.A1(net2121),
    .A2(_1779_),
    .B1(net2083),
    .Y(_1780_));
 sky130_fd_sc_hd__mux2_1 _4138_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[3] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[3] ),
    .S(net376),
    .X(_1781_));
 sky130_fd_sc_hd__nor2_1 _4139_ (.A(net2154),
    .B(_1781_),
    .Y(_1782_));
 sky130_fd_sc_hd__and2_1 _4140_ (.A(net2154),
    .B(_1781_),
    .X(_1783_));
 sky130_fd_sc_hd__or2_1 _4141_ (.A(net2155),
    .B(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__mux2_1 _4142_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[2] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[2] ),
    .S(net375),
    .X(_1785_));
 sky130_fd_sc_hd__and2_2 _4143_ (.A(net2169),
    .B(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__and3_1 _4144_ (.A(net2136),
    .B(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ),
    .C(net375),
    .X(_1787_));
 sky130_fd_sc_hd__a21oi_1 _4145_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ),
    .A2(net375),
    .B1(net2136),
    .Y(_1788_));
 sky130_fd_sc_hd__or2_1 _4146_ (.A(_1787_),
    .B(net2137),
    .X(_1789_));
 sky130_fd_sc_hd__nand3_1 _4147_ (.A(net1878),
    .B(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ),
    .C(net375),
    .Y(_1790_));
 sky130_fd_sc_hd__nor2_1 _4148_ (.A(_1789_),
    .B(_1790_),
    .Y(_1791_));
 sky130_fd_sc_hd__or2_1 _4149_ (.A(_1787_),
    .B(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__nor2_1 _4150_ (.A(net2169),
    .B(_1785_),
    .Y(_1793_));
 sky130_fd_sc_hd__or2_1 _4151_ (.A(_1786_),
    .B(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__and2b_2 _4152_ (.A_N(_1794_),
    .B(_1792_),
    .X(_1795_));
 sky130_fd_sc_hd__or2_1 _4153_ (.A(_1786_),
    .B(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__o21ba_1 _4154_ (.A1(_1786_),
    .A2(_1795_),
    .B1_N(_1784_),
    .X(_1797_));
 sky130_fd_sc_hd__xnor2_1 _4155_ (.A(net2156),
    .B(_1796_),
    .Y(_1798_));
 sky130_fd_sc_hd__mux2_1 _4156_ (.A0(_1798_),
    .A1(net2004),
    .S(net179),
    .X(_1799_));
 sky130_fd_sc_hd__and2b_1 _4157_ (.A_N(_1792_),
    .B(_1794_),
    .X(_1800_));
 sky130_fd_sc_hd__nor2_4 _4158_ (.A(_1795_),
    .B(_1800_),
    .Y(_1801_));
 sky130_fd_sc_hd__mux2_8 _4159_ (.A0(_1801_),
    .A1(net2100),
    .S(net174),
    .X(_1802_));
 sky130_fd_sc_hd__inv_2 _4160_ (.A(_1802_),
    .Y(_1803_));
 sky130_fd_sc_hd__nand2_1 _4161_ (.A(_1799_),
    .B(_1802_),
    .Y(_1804_));
 sky130_fd_sc_hd__mux2_1 _4162_ (.A0(net2258),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[4] ),
    .S(net375),
    .X(_1805_));
 sky130_fd_sc_hd__nor2_1 _4163_ (.A(net2229),
    .B(_1805_),
    .Y(_1806_));
 sky130_fd_sc_hd__and2_1 _4164_ (.A(net2229),
    .B(net2259),
    .X(_1807_));
 sky130_fd_sc_hd__or2_1 _4165_ (.A(_1806_),
    .B(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__o21ba_1 _4166_ (.A1(_1783_),
    .A2(_1797_),
    .B1_N(_1808_),
    .X(_1809_));
 sky130_fd_sc_hd__or3b_1 _4167_ (.A(_1783_),
    .B(_1797_),
    .C_N(_1808_),
    .X(_1810_));
 sky130_fd_sc_hd__and2b_1 _4168_ (.A_N(_1809_),
    .B(_1810_),
    .X(_1811_));
 sky130_fd_sc_hd__mux2_1 _4169_ (.A0(_1811_),
    .A1(net2054),
    .S(net179),
    .X(_1812_));
 sky130_fd_sc_hd__nand2b_2 _4170_ (.A_N(_1804_),
    .B(_1812_),
    .Y(_1813_));
 sky130_fd_sc_hd__mux2_1 _4171_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[5] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[5] ),
    .S(net375),
    .X(_1814_));
 sky130_fd_sc_hd__nor2_1 _4172_ (.A(net2170),
    .B(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__and2_1 _4173_ (.A(net2170),
    .B(_1814_),
    .X(_1816_));
 sky130_fd_sc_hd__or2_1 _4174_ (.A(_1815_),
    .B(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__o21ba_1 _4175_ (.A1(_1807_),
    .A2(_1809_),
    .B1_N(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__or3b_1 _4176_ (.A(_1807_),
    .B(_1809_),
    .C_N(_1817_),
    .X(_1819_));
 sky130_fd_sc_hd__and2b_1 _4177_ (.A_N(_1818_),
    .B(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__mux2_2 _4178_ (.A0(_1820_),
    .A1(net1993),
    .S(net176),
    .X(_1821_));
 sky130_fd_sc_hd__inv_2 _4179_ (.A(_1821_),
    .Y(_1822_));
 sky130_fd_sc_hd__mux2_1 _4180_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[6] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ),
    .S(net376),
    .X(_1823_));
 sky130_fd_sc_hd__nor2_1 _4181_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ),
    .B(_1823_),
    .Y(_1824_));
 sky130_fd_sc_hd__and2_1 _4182_ (.A(net2175),
    .B(_1823_),
    .X(_1825_));
 sky130_fd_sc_hd__or2_1 _4183_ (.A(_1824_),
    .B(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__o21ba_1 _4184_ (.A1(_1816_),
    .A2(_1818_),
    .B1_N(_1826_),
    .X(_1827_));
 sky130_fd_sc_hd__or3b_1 _4185_ (.A(net2171),
    .B(_1818_),
    .C_N(_1826_),
    .X(_1828_));
 sky130_fd_sc_hd__and2b_1 _4186_ (.A_N(_1827_),
    .B(net2172),
    .X(_1829_));
 sky130_fd_sc_hd__mux2_1 _4187_ (.A0(_1829_),
    .A1(net1992),
    .S(net178),
    .X(_1830_));
 sky130_fd_sc_hd__inv_2 _4188_ (.A(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__or3_1 _4189_ (.A(_1813_),
    .B(_1822_),
    .C(_1831_),
    .X(_1832_));
 sky130_fd_sc_hd__mux2_1 _4190_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[7] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[7] ),
    .S(\U_DATAPATH.U_ID_EX.o_addr_src_EX ),
    .X(_1833_));
 sky130_fd_sc_hd__nor2_1 _4191_ (.A(net2160),
    .B(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__and2_1 _4192_ (.A(net2160),
    .B(_1833_),
    .X(_1835_));
 sky130_fd_sc_hd__or2_1 _4193_ (.A(_1834_),
    .B(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__o21ba_1 _4194_ (.A1(_1825_),
    .A2(_1827_),
    .B1_N(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__or3b_1 _4195_ (.A(net2176),
    .B(_1827_),
    .C_N(_1836_),
    .X(_1838_));
 sky130_fd_sc_hd__and2b_1 _4196_ (.A_N(_1837_),
    .B(_1838_),
    .X(_1839_));
 sky130_fd_sc_hd__mux2_1 _4197_ (.A0(_1839_),
    .A1(net2017),
    .S(net179),
    .X(_1840_));
 sky130_fd_sc_hd__nand2b_1 _4198_ (.A_N(_1832_),
    .B(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__mux2_1 _4199_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[8] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[8] ),
    .S(net376),
    .X(_1842_));
 sky130_fd_sc_hd__nor2_1 _4200_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ),
    .B(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__and2_1 _4201_ (.A(net2224),
    .B(_1842_),
    .X(_1844_));
 sky130_fd_sc_hd__or2_1 _4202_ (.A(_1843_),
    .B(_1844_),
    .X(_1845_));
 sky130_fd_sc_hd__o21ba_1 _4203_ (.A1(net2161),
    .A2(_1837_),
    .B1_N(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__or3b_1 _4204_ (.A(net2161),
    .B(_1837_),
    .C_N(_1845_),
    .X(_1847_));
 sky130_fd_sc_hd__nand2b_1 _4205_ (.A_N(_1846_),
    .B(net2162),
    .Y(_1848_));
 sky130_fd_sc_hd__inv_2 _4206_ (.A(_1848_),
    .Y(_1849_));
 sky130_fd_sc_hd__mux2_1 _4207_ (.A0(_1849_),
    .A1(net2061),
    .S(net179),
    .X(_1850_));
 sky130_fd_sc_hd__nand2b_1 _4208_ (.A_N(_1841_),
    .B(_1850_),
    .Y(_1851_));
 sky130_fd_sc_hd__mux2_1 _4209_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[9] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ),
    .S(net375),
    .X(_1852_));
 sky130_fd_sc_hd__nor2_1 _4210_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ),
    .B(_1852_),
    .Y(_1853_));
 sky130_fd_sc_hd__and2_1 _4211_ (.A(net2240),
    .B(_1852_),
    .X(_1854_));
 sky130_fd_sc_hd__or2_1 _4212_ (.A(_1853_),
    .B(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__o21ba_1 _4213_ (.A1(_1844_),
    .A2(_1846_),
    .B1_N(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__or3b_1 _4214_ (.A(net2225),
    .B(_1846_),
    .C_N(_1855_),
    .X(_1857_));
 sky130_fd_sc_hd__and2b_1 _4215_ (.A_N(_1856_),
    .B(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__mux2_1 _4216_ (.A0(_1858_),
    .A1(net2013),
    .S(net180),
    .X(_1859_));
 sky130_fd_sc_hd__and2b_1 _4217_ (.A_N(_1851_),
    .B(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__mux2_1 _4218_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[10] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[10] ),
    .S(\U_DATAPATH.U_ID_EX.o_addr_src_EX ),
    .X(_1861_));
 sky130_fd_sc_hd__nor2_1 _4219_ (.A(net2189),
    .B(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__and2_1 _4220_ (.A(net2189),
    .B(_1861_),
    .X(_1863_));
 sky130_fd_sc_hd__or2_1 _4221_ (.A(_1862_),
    .B(_1863_),
    .X(_1864_));
 sky130_fd_sc_hd__o21ba_1 _4222_ (.A1(_1854_),
    .A2(_1856_),
    .B1_N(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__or3b_1 _4223_ (.A(net2241),
    .B(_1856_),
    .C_N(_1864_),
    .X(_1866_));
 sky130_fd_sc_hd__and2b_1 _4224_ (.A_N(_1865_),
    .B(_1866_),
    .X(_1867_));
 sky130_fd_sc_hd__mux2_1 _4225_ (.A0(_1867_),
    .A1(net2044),
    .S(net176),
    .X(_1868_));
 sky130_fd_sc_hd__and2_1 _4226_ (.A(_1860_),
    .B(_1868_),
    .X(_1869_));
 sky130_fd_sc_hd__mux2_1 _4227_ (.A0(net2348),
    .A1(net2341),
    .S(\U_DATAPATH.U_ID_EX.o_addr_src_EX ),
    .X(_1870_));
 sky130_fd_sc_hd__nor2_1 _4228_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ),
    .B(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__and2_1 _4229_ (.A(net2214),
    .B(_1870_),
    .X(_1872_));
 sky130_fd_sc_hd__or2_1 _4230_ (.A(_1871_),
    .B(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__o21ba_1 _4231_ (.A1(_1863_),
    .A2(_1865_),
    .B1_N(_1873_),
    .X(_1874_));
 sky130_fd_sc_hd__or3b_1 _4232_ (.A(net2190),
    .B(_1865_),
    .C_N(_1873_),
    .X(_1875_));
 sky130_fd_sc_hd__and2b_1 _4233_ (.A_N(_1874_),
    .B(net2191),
    .X(_1876_));
 sky130_fd_sc_hd__mux2_1 _4234_ (.A0(_1876_),
    .A1(net2060),
    .S(net175),
    .X(_1877_));
 sky130_fd_sc_hd__nand2_1 _4235_ (.A(_1869_),
    .B(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__mux2_1 _4236_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[12] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ),
    .S(net375),
    .X(_1879_));
 sky130_fd_sc_hd__nor2_1 _4237_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ),
    .B(_1879_),
    .Y(_1880_));
 sky130_fd_sc_hd__and2_1 _4238_ (.A(net2164),
    .B(_1879_),
    .X(_1881_));
 sky130_fd_sc_hd__or2_1 _4239_ (.A(_1880_),
    .B(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__o21ba_1 _4240_ (.A1(_1872_),
    .A2(_1874_),
    .B1_N(_1882_),
    .X(_1883_));
 sky130_fd_sc_hd__or3b_1 _4241_ (.A(_1872_),
    .B(_1874_),
    .C_N(_1882_),
    .X(_1884_));
 sky130_fd_sc_hd__and2b_1 _4242_ (.A_N(_1883_),
    .B(_1884_),
    .X(_1885_));
 sky130_fd_sc_hd__mux2_2 _4243_ (.A0(_1885_),
    .A1(net2027),
    .S(net179),
    .X(_1886_));
 sky130_fd_sc_hd__mux2_1 _4244_ (.A0(net2237),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ),
    .S(net375),
    .X(_1887_));
 sky130_fd_sc_hd__nor2_1 _4245_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ),
    .B(_1887_),
    .Y(_1888_));
 sky130_fd_sc_hd__and2_1 _4246_ (.A(net2199),
    .B(net2238),
    .X(_1889_));
 sky130_fd_sc_hd__or2_1 _4247_ (.A(_1888_),
    .B(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__o21ba_1 _4248_ (.A1(_1881_),
    .A2(_1883_),
    .B1_N(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__or3b_1 _4249_ (.A(net2165),
    .B(_1883_),
    .C_N(_1890_),
    .X(_1892_));
 sky130_fd_sc_hd__and2b_1 _4250_ (.A_N(_1891_),
    .B(net2166),
    .X(_1893_));
 sky130_fd_sc_hd__mux2_2 _4251_ (.A0(_1893_),
    .A1(net1971),
    .S(net175),
    .X(_1894_));
 sky130_fd_sc_hd__nand3b_1 _4252_ (.A_N(_1878_),
    .B(_1886_),
    .C(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__mux2_1 _4253_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[14] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[14] ),
    .S(net375),
    .X(_1896_));
 sky130_fd_sc_hd__nor2_1 _4254_ (.A(net2193),
    .B(_1896_),
    .Y(_1897_));
 sky130_fd_sc_hd__and2_1 _4255_ (.A(net2193),
    .B(_1896_),
    .X(_1898_));
 sky130_fd_sc_hd__or2_1 _4256_ (.A(_1897_),
    .B(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__o21ba_1 _4257_ (.A1(_1889_),
    .A2(_1891_),
    .B1_N(_1899_),
    .X(_1900_));
 sky130_fd_sc_hd__or3b_1 _4258_ (.A(_1889_),
    .B(_1891_),
    .C_N(_1899_),
    .X(_1901_));
 sky130_fd_sc_hd__nand2b_1 _4259_ (.A_N(_1900_),
    .B(net2239),
    .Y(_1902_));
 sky130_fd_sc_hd__inv_2 _4260_ (.A(_1902_),
    .Y(_1903_));
 sky130_fd_sc_hd__mux2_1 _4261_ (.A0(_1903_),
    .A1(net1989),
    .S(net175),
    .X(_1904_));
 sky130_fd_sc_hd__and2b_1 _4262_ (.A_N(_1895_),
    .B(_1904_),
    .X(_1905_));
 sky130_fd_sc_hd__mux2_1 _4263_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[15] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[15] ),
    .S(net375),
    .X(_1906_));
 sky130_fd_sc_hd__nor2_1 _4264_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ),
    .B(_1906_),
    .Y(_1907_));
 sky130_fd_sc_hd__and2_1 _4265_ (.A(net2226),
    .B(_1906_),
    .X(_1908_));
 sky130_fd_sc_hd__or2_1 _4266_ (.A(_1907_),
    .B(_1908_),
    .X(_1909_));
 sky130_fd_sc_hd__o21ba_1 _4267_ (.A1(_1898_),
    .A2(_1900_),
    .B1_N(_1909_),
    .X(_1910_));
 sky130_fd_sc_hd__or3b_1 _4268_ (.A(net2194),
    .B(_1900_),
    .C_N(_1909_),
    .X(_1911_));
 sky130_fd_sc_hd__and2b_1 _4269_ (.A_N(_1910_),
    .B(net2195),
    .X(_1912_));
 sky130_fd_sc_hd__mux2_2 _4270_ (.A0(_1912_),
    .A1(net2015),
    .S(net175),
    .X(_1913_));
 sky130_fd_sc_hd__and2_2 _4271_ (.A(_1905_),
    .B(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__mux2_1 _4272_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[16] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ),
    .S(net375),
    .X(_1915_));
 sky130_fd_sc_hd__nor2_1 _4273_ (.A(net2075),
    .B(_1915_),
    .Y(_1916_));
 sky130_fd_sc_hd__and2_1 _4274_ (.A(net2075),
    .B(_1915_),
    .X(_1917_));
 sky130_fd_sc_hd__or2_1 _4275_ (.A(_1916_),
    .B(_1917_),
    .X(_1918_));
 sky130_fd_sc_hd__o21ba_1 _4276_ (.A1(_1908_),
    .A2(_1910_),
    .B1_N(_1918_),
    .X(_1919_));
 sky130_fd_sc_hd__or3b_1 _4277_ (.A(net2227),
    .B(_1910_),
    .C_N(_1918_),
    .X(_1920_));
 sky130_fd_sc_hd__and2b_1 _4278_ (.A_N(_1919_),
    .B(net2228),
    .X(_1921_));
 sky130_fd_sc_hd__mux2_2 _4279_ (.A0(_1921_),
    .A1(net2023),
    .S(net177),
    .X(_1922_));
 sky130_fd_sc_hd__mux2_1 _4280_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[17] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ),
    .S(net375),
    .X(_1923_));
 sky130_fd_sc_hd__nor2_1 _4281_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ),
    .B(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__and2_1 _4282_ (.A(net2200),
    .B(_1923_),
    .X(_1925_));
 sky130_fd_sc_hd__or2_1 _4283_ (.A(_1924_),
    .B(_1925_),
    .X(_1926_));
 sky130_fd_sc_hd__o21ba_1 _4284_ (.A1(net2076),
    .A2(_1919_),
    .B1_N(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__or3b_1 _4285_ (.A(net2076),
    .B(_1919_),
    .C_N(_1926_),
    .X(_1928_));
 sky130_fd_sc_hd__nand2b_1 _4286_ (.A_N(_1927_),
    .B(net2077),
    .Y(_1929_));
 sky130_fd_sc_hd__inv_2 _4287_ (.A(_1929_),
    .Y(_1930_));
 sky130_fd_sc_hd__mux2_1 _4288_ (.A0(_1930_),
    .A1(net2068),
    .S(net178),
    .X(_1931_));
 sky130_fd_sc_hd__and3_1 _4289_ (.A(_1914_),
    .B(_1922_),
    .C(_1931_),
    .X(_1932_));
 sky130_fd_sc_hd__mux2_1 _4290_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[18] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[18] ),
    .S(net375),
    .X(_1933_));
 sky130_fd_sc_hd__nor2_1 _4291_ (.A(net2148),
    .B(_1933_),
    .Y(_1934_));
 sky130_fd_sc_hd__and2_1 _4292_ (.A(net2148),
    .B(_1933_),
    .X(_1935_));
 sky130_fd_sc_hd__or2_1 _4293_ (.A(_1934_),
    .B(_1935_),
    .X(_1936_));
 sky130_fd_sc_hd__o21ba_1 _4294_ (.A1(_1925_),
    .A2(_1927_),
    .B1_N(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__or3b_1 _4295_ (.A(net2201),
    .B(_1927_),
    .C_N(_1936_),
    .X(_1938_));
 sky130_fd_sc_hd__and2b_1 _4296_ (.A_N(_1937_),
    .B(_1938_),
    .X(_1939_));
 sky130_fd_sc_hd__mux2_4 _4297_ (.A0(_1939_),
    .A1(net2070),
    .S(net178),
    .X(_1940_));
 sky130_fd_sc_hd__and2_4 _4298_ (.A(_1932_),
    .B(_1940_),
    .X(_1941_));
 sky130_fd_sc_hd__mux2_1 _4299_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[19] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[19] ),
    .S(net375),
    .X(_1942_));
 sky130_fd_sc_hd__nor2_1 _4300_ (.A(net2132),
    .B(_1942_),
    .Y(_1943_));
 sky130_fd_sc_hd__and2_1 _4301_ (.A(net2132),
    .B(_1942_),
    .X(_1944_));
 sky130_fd_sc_hd__or2_1 _4302_ (.A(_1943_),
    .B(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__o21ba_2 _4303_ (.A1(_1935_),
    .A2(_1937_),
    .B1_N(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__or3b_1 _4304_ (.A(net2149),
    .B(_1937_),
    .C_N(_1945_),
    .X(_1947_));
 sky130_fd_sc_hd__and2b_1 _4305_ (.A_N(_1946_),
    .B(net2150),
    .X(_1948_));
 sky130_fd_sc_hd__mux2_1 _4306_ (.A0(_1948_),
    .A1(net2024),
    .S(net177),
    .X(_1949_));
 sky130_fd_sc_hd__nand2_1 _4307_ (.A(_1941_),
    .B(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__mux2_1 _4308_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[20] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[20] ),
    .S(net376),
    .X(_1951_));
 sky130_fd_sc_hd__nor2_1 _4309_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ),
    .B(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__and2_1 _4310_ (.A(net2243),
    .B(_1951_),
    .X(_1953_));
 sky130_fd_sc_hd__or2_1 _4311_ (.A(_1952_),
    .B(_1953_),
    .X(_1954_));
 sky130_fd_sc_hd__o21ba_1 _4312_ (.A1(net2133),
    .A2(_1946_),
    .B1_N(_1954_),
    .X(_1955_));
 sky130_fd_sc_hd__or3b_1 _4313_ (.A(net2133),
    .B(_1946_),
    .C_N(_1954_),
    .X(_1956_));
 sky130_fd_sc_hd__nand2b_1 _4314_ (.A_N(_1955_),
    .B(net2134),
    .Y(_1957_));
 sky130_fd_sc_hd__inv_2 _4315_ (.A(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__mux2_4 _4316_ (.A0(_1958_),
    .A1(net2064),
    .S(net183),
    .X(_1959_));
 sky130_fd_sc_hd__and3_4 _4317_ (.A(_1941_),
    .B(_1949_),
    .C(_1959_),
    .X(_1960_));
 sky130_fd_sc_hd__mux2_1 _4318_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[21] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[21] ),
    .S(net376),
    .X(_1961_));
 sky130_fd_sc_hd__nor2_1 _4319_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ),
    .B(_1961_),
    .Y(_1962_));
 sky130_fd_sc_hd__and2_1 _4320_ (.A(net2263),
    .B(_1961_),
    .X(_1963_));
 sky130_fd_sc_hd__or2_1 _4321_ (.A(_1962_),
    .B(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__o21ba_1 _4322_ (.A1(net2244),
    .A2(_1955_),
    .B1_N(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__or3b_1 _4323_ (.A(net2244),
    .B(_1955_),
    .C_N(_1964_),
    .X(_1966_));
 sky130_fd_sc_hd__and2b_1 _4324_ (.A_N(_1965_),
    .B(net2245),
    .X(_1967_));
 sky130_fd_sc_hd__mux2_1 _4325_ (.A0(_1967_),
    .A1(net1874),
    .S(net172),
    .X(_1968_));
 sky130_fd_sc_hd__and2_1 _4326_ (.A(_1960_),
    .B(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__mux2_1 _4327_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[22] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ),
    .S(net376),
    .X(_1970_));
 sky130_fd_sc_hd__nor2_1 _4328_ (.A(net2181),
    .B(_1970_),
    .Y(_1971_));
 sky130_fd_sc_hd__and2_1 _4329_ (.A(net2181),
    .B(_1970_),
    .X(_1972_));
 sky130_fd_sc_hd__or2_1 _4330_ (.A(_1971_),
    .B(net2182),
    .X(_1973_));
 sky130_fd_sc_hd__o21ba_1 _4331_ (.A1(net2264),
    .A2(_1965_),
    .B1_N(_1973_),
    .X(_1974_));
 sky130_fd_sc_hd__or3b_1 _4332_ (.A(net2264),
    .B(_1965_),
    .C_N(_1973_),
    .X(_1975_));
 sky130_fd_sc_hd__nand2b_1 _4333_ (.A_N(_1974_),
    .B(net2265),
    .Y(_1976_));
 sky130_fd_sc_hd__inv_2 _4334_ (.A(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hd__mux2_1 _4335_ (.A0(_1977_),
    .A1(net1988),
    .S(net172),
    .X(_1978_));
 sky130_fd_sc_hd__mux2_1 _4336_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[23] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[23] ),
    .S(net376),
    .X(_1979_));
 sky130_fd_sc_hd__nor2_1 _4337_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ),
    .B(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__and2_1 _4338_ (.A(net2210),
    .B(_1979_),
    .X(_1981_));
 sky130_fd_sc_hd__or2_1 _4339_ (.A(_1980_),
    .B(_1981_),
    .X(_1982_));
 sky130_fd_sc_hd__o21ba_1 _4340_ (.A1(_1972_),
    .A2(_1974_),
    .B1_N(_1982_),
    .X(_1983_));
 sky130_fd_sc_hd__or3b_1 _4341_ (.A(net2182),
    .B(_1974_),
    .C_N(_1982_),
    .X(_1984_));
 sky130_fd_sc_hd__and2b_1 _4342_ (.A_N(_1983_),
    .B(net2183),
    .X(_1985_));
 sky130_fd_sc_hd__mux2_2 _4343_ (.A0(_1985_),
    .A1(net2021),
    .S(net172),
    .X(_1986_));
 sky130_fd_sc_hd__and3_1 _4344_ (.A(_1969_),
    .B(_1978_),
    .C(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__mux2_1 _4345_ (.A0(net2334),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ),
    .S(net376),
    .X(_1988_));
 sky130_fd_sc_hd__nor2_1 _4346_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ),
    .B(_1988_),
    .Y(_1989_));
 sky130_fd_sc_hd__and2_1 _4347_ (.A(net2301),
    .B(_1988_),
    .X(_1990_));
 sky130_fd_sc_hd__or2_1 _4348_ (.A(_1989_),
    .B(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__o21ba_1 _4349_ (.A1(_1981_),
    .A2(_1983_),
    .B1_N(_1991_),
    .X(_1992_));
 sky130_fd_sc_hd__or3b_1 _4350_ (.A(net2211),
    .B(_1983_),
    .C_N(_1991_),
    .X(_1993_));
 sky130_fd_sc_hd__and2b_1 _4351_ (.A_N(_1992_),
    .B(net2212),
    .X(_1994_));
 sky130_fd_sc_hd__mux2_1 _4352_ (.A0(_1994_),
    .A1(net2059),
    .S(net172),
    .X(_1995_));
 sky130_fd_sc_hd__and2_1 _4353_ (.A(_1987_),
    .B(_1995_),
    .X(_1996_));
 sky130_fd_sc_hd__mux2_1 _4354_ (.A0(net2318),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[25] ),
    .S(net376),
    .X(_1997_));
 sky130_fd_sc_hd__nor2_1 _4355_ (.A(net2281),
    .B(_1997_),
    .Y(_1998_));
 sky130_fd_sc_hd__and2_1 _4356_ (.A(net2281),
    .B(net2319),
    .X(_1999_));
 sky130_fd_sc_hd__or2_1 _4357_ (.A(_1998_),
    .B(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__o21ba_1 _4358_ (.A1(_1990_),
    .A2(_1992_),
    .B1_N(_2000_),
    .X(_2001_));
 sky130_fd_sc_hd__or3b_1 _4359_ (.A(_1990_),
    .B(_1992_),
    .C_N(_2000_),
    .X(_2002_));
 sky130_fd_sc_hd__and2b_1 _4360_ (.A_N(_2001_),
    .B(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__mux2_1 _4361_ (.A0(_2003_),
    .A1(net2055),
    .S(net171),
    .X(_2004_));
 sky130_fd_sc_hd__and3_1 _4362_ (.A(_1987_),
    .B(_1995_),
    .C(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__mux2_1 _4363_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[26] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[26] ),
    .S(net376),
    .X(_2006_));
 sky130_fd_sc_hd__nor2_1 _4364_ (.A(net2233),
    .B(_2006_),
    .Y(_2007_));
 sky130_fd_sc_hd__and2_1 _4365_ (.A(net2233),
    .B(_2006_),
    .X(_2008_));
 sky130_fd_sc_hd__or2_1 _4366_ (.A(_2007_),
    .B(_2008_),
    .X(_2009_));
 sky130_fd_sc_hd__o21ba_1 _4367_ (.A1(_1999_),
    .A2(_2001_),
    .B1_N(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__or3b_1 _4368_ (.A(_1999_),
    .B(_2001_),
    .C_N(_2009_),
    .X(_2011_));
 sky130_fd_sc_hd__and2b_1 _4369_ (.A_N(_2010_),
    .B(_2011_),
    .X(_2012_));
 sky130_fd_sc_hd__mux2_1 _4370_ (.A0(_2012_),
    .A1(net2052),
    .S(net173),
    .X(_2013_));
 sky130_fd_sc_hd__and2_1 _4371_ (.A(_2005_),
    .B(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__mux2_1 _4372_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[27] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[27] ),
    .S(net376),
    .X(_2015_));
 sky130_fd_sc_hd__nor2_1 _4373_ (.A(net2186),
    .B(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__and2_1 _4374_ (.A(net2186),
    .B(_2015_),
    .X(_2017_));
 sky130_fd_sc_hd__or2_1 _4375_ (.A(_2016_),
    .B(_2017_),
    .X(_2018_));
 sky130_fd_sc_hd__o21ba_1 _4376_ (.A1(_2008_),
    .A2(_2010_),
    .B1_N(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__or3b_1 _4377_ (.A(net2234),
    .B(_2010_),
    .C_N(_2018_),
    .X(_2020_));
 sky130_fd_sc_hd__and2b_1 _4378_ (.A_N(_2019_),
    .B(net2235),
    .X(_2021_));
 sky130_fd_sc_hd__mux2_1 _4379_ (.A0(_2021_),
    .A1(net2029),
    .S(net173),
    .X(_2022_));
 sky130_fd_sc_hd__and3_1 _4380_ (.A(_2005_),
    .B(_2013_),
    .C(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__mux2_1 _4381_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[28] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[28] ),
    .S(net376),
    .X(_2024_));
 sky130_fd_sc_hd__nor2_1 _4382_ (.A(net2040),
    .B(_2024_),
    .Y(_2025_));
 sky130_fd_sc_hd__and2_1 _4383_ (.A(net2040),
    .B(_2024_),
    .X(_2026_));
 sky130_fd_sc_hd__or2_1 _4384_ (.A(_2025_),
    .B(_2026_),
    .X(_2027_));
 sky130_fd_sc_hd__o21ba_1 _4385_ (.A1(_2017_),
    .A2(_2019_),
    .B1_N(_2027_),
    .X(_2028_));
 sky130_fd_sc_hd__or3b_1 _4386_ (.A(net2187),
    .B(_2019_),
    .C_N(_2027_),
    .X(_2029_));
 sky130_fd_sc_hd__and2b_1 _4387_ (.A_N(_2028_),
    .B(net2188),
    .X(_2030_));
 sky130_fd_sc_hd__mux2_1 _4388_ (.A0(_2030_),
    .A1(net1954),
    .S(net171),
    .X(_2031_));
 sky130_fd_sc_hd__and2_1 _4389_ (.A(_2023_),
    .B(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__mux2_1 _4390_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[29] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[29] ),
    .S(net376),
    .X(_2033_));
 sky130_fd_sc_hd__nor2_1 _4391_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ),
    .B(_2033_),
    .Y(_2034_));
 sky130_fd_sc_hd__and2_1 _4392_ (.A(net2216),
    .B(_2033_),
    .X(_2035_));
 sky130_fd_sc_hd__or2_1 _4393_ (.A(_2034_),
    .B(_2035_),
    .X(_2036_));
 sky130_fd_sc_hd__o21ba_1 _4394_ (.A1(_2026_),
    .A2(_2028_),
    .B1_N(_2036_),
    .X(_2037_));
 sky130_fd_sc_hd__or3b_1 _4395_ (.A(net2041),
    .B(_2028_),
    .C_N(_2036_),
    .X(_2038_));
 sky130_fd_sc_hd__and2b_1 _4396_ (.A_N(_2037_),
    .B(net2042),
    .X(_2039_));
 sky130_fd_sc_hd__mux2_1 _4397_ (.A0(_2039_),
    .A1(net2031),
    .S(net171),
    .X(_2040_));
 sky130_fd_sc_hd__and3_1 _4398_ (.A(_2023_),
    .B(_2031_),
    .C(_2040_),
    .X(_2041_));
 sky130_fd_sc_hd__mux2_1 _4399_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[30] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ),
    .S(net376),
    .X(_2042_));
 sky130_fd_sc_hd__xnor2_1 _4400_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ),
    .B(_2042_),
    .Y(_2043_));
 sky130_fd_sc_hd__o21ba_1 _4401_ (.A1(_2035_),
    .A2(_2037_),
    .B1_N(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__or3b_1 _4402_ (.A(net2217),
    .B(_2037_),
    .C_N(_2043_),
    .X(_2045_));
 sky130_fd_sc_hd__and2b_1 _4403_ (.A_N(_2044_),
    .B(net2218),
    .X(_2046_));
 sky130_fd_sc_hd__mux2_1 _4404_ (.A0(_2046_),
    .A1(net1887),
    .S(net171),
    .X(_2047_));
 sky130_fd_sc_hd__and2_1 _4405_ (.A(_2041_),
    .B(_2047_),
    .X(_2048_));
 sky130_fd_sc_hd__a21o_1 _4406_ (.A1(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ),
    .A2(_2042_),
    .B1(_2044_),
    .X(_2049_));
 sky130_fd_sc_hd__xnor2_1 _4407_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ),
    .B(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__mux2_1 _4408_ (.A0(net2247),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ),
    .S(net376),
    .X(_2051_));
 sky130_fd_sc_hd__xnor2_1 _4409_ (.A(_2050_),
    .B(net2248),
    .Y(_2052_));
 sky130_fd_sc_hd__mux2_1 _4410_ (.A0(net2249),
    .A1(net2036),
    .S(net171),
    .X(_2053_));
 sky130_fd_sc_hd__or2_1 _4411_ (.A(net390),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .X(_2054_));
 sky130_fd_sc_hd__nand2_1 _4412_ (.A(net390),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .Y(_2055_));
 sky130_fd_sc_hd__or2_1 _4413_ (.A(net402),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .X(_2056_));
 sky130_fd_sc_hd__nand2_1 _4414_ (.A(net402),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .Y(_2057_));
 sky130_fd_sc_hd__a22o_1 _4415_ (.A1(_2054_),
    .A2(_2055_),
    .B1(_2056_),
    .B2(_2057_),
    .X(_2058_));
 sky130_fd_sc_hd__or2_1 _4416_ (.A(net379),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .X(_2059_));
 sky130_fd_sc_hd__nand2_1 _4417_ (.A(net379),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .Y(_2060_));
 sky130_fd_sc_hd__or2_1 _4418_ (.A(net383),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .X(_2061_));
 sky130_fd_sc_hd__nand2_1 _4419_ (.A(net383),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .Y(_2062_));
 sky130_fd_sc_hd__a22o_1 _4420_ (.A1(_2059_),
    .A2(_2060_),
    .B1(_2061_),
    .B2(_2062_),
    .X(_2063_));
 sky130_fd_sc_hd__or2_1 _4421_ (.A(net429),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .X(_2064_));
 sky130_fd_sc_hd__nand2_1 _4422_ (.A(net429),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .Y(_2065_));
 sky130_fd_sc_hd__or2_1 _4423_ (.A(net407),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .X(_2066_));
 sky130_fd_sc_hd__nand2_1 _4424_ (.A(net407),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .Y(_2067_));
 sky130_fd_sc_hd__or2_1 _4425_ (.A(net420),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .X(_2068_));
 sky130_fd_sc_hd__nand2_1 _4426_ (.A(net420),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .Y(_2069_));
 sky130_fd_sc_hd__or2_1 _4427_ (.A(net411),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .X(_2070_));
 sky130_fd_sc_hd__nand2_1 _4428_ (.A(net411),
    .B(net2074),
    .Y(_2071_));
 sky130_fd_sc_hd__a22o_1 _4429_ (.A1(_2064_),
    .A2(_2065_),
    .B1(_2068_),
    .B2(_2069_),
    .X(_2072_));
 sky130_fd_sc_hd__a22o_1 _4430_ (.A1(_2066_),
    .A2(_2067_),
    .B1(_2070_),
    .B2(_2071_),
    .X(_2073_));
 sky130_fd_sc_hd__o22a_2 _4431_ (.A1(_2058_),
    .A2(_2063_),
    .B1(_2072_),
    .B2(_2073_),
    .X(_2074_));
 sky130_fd_sc_hd__nor3b_4 _4432_ (.A(net610),
    .B(_2074_),
    .C_N(net1987),
    .Y(_2075_));
 sky130_fd_sc_hd__or3b_1 _4433_ (.A(net610),
    .B(_2074_),
    .C_N(net1987),
    .X(_2076_));
 sky130_fd_sc_hd__nor2_1 _4434_ (.A(_2048_),
    .B(net292),
    .Y(_2077_));
 sky130_fd_sc_hd__nand2_1 _4435_ (.A(_2048_),
    .B(_2053_),
    .Y(_2078_));
 sky130_fd_sc_hd__o21a_1 _4436_ (.A1(_2048_),
    .A2(_2053_),
    .B1(net271),
    .X(_2079_));
 sky130_fd_sc_hd__a22o_1 _4437_ (.A1(net2036),
    .A2(net292),
    .B1(_2078_),
    .B2(_2079_),
    .X(_1143_));
 sky130_fd_sc_hd__or2_1 _4438_ (.A(_2041_),
    .B(_2047_),
    .X(_2080_));
 sky130_fd_sc_hd__a22o_1 _4439_ (.A1(net1887),
    .A2(net292),
    .B1(_2077_),
    .B2(_2080_),
    .X(_1142_));
 sky130_fd_sc_hd__or2_1 _4440_ (.A(_2032_),
    .B(_2040_),
    .X(_2081_));
 sky130_fd_sc_hd__nor2_1 _4441_ (.A(_2041_),
    .B(net292),
    .Y(_2082_));
 sky130_fd_sc_hd__a22o_1 _4442_ (.A1(net2031),
    .A2(net292),
    .B1(_2081_),
    .B2(_2082_),
    .X(_1141_));
 sky130_fd_sc_hd__or2_1 _4443_ (.A(_2023_),
    .B(_2031_),
    .X(_2083_));
 sky130_fd_sc_hd__nor2_1 _4444_ (.A(_2032_),
    .B(net292),
    .Y(_2084_));
 sky130_fd_sc_hd__a22o_1 _4445_ (.A1(net1954),
    .A2(net292),
    .B1(_2083_),
    .B2(_2084_),
    .X(_1140_));
 sky130_fd_sc_hd__or2_1 _4446_ (.A(_2014_),
    .B(_2022_),
    .X(_2085_));
 sky130_fd_sc_hd__nor2_1 _4447_ (.A(_2023_),
    .B(net293),
    .Y(_2086_));
 sky130_fd_sc_hd__a22o_1 _4448_ (.A1(net2029),
    .A2(net293),
    .B1(_2085_),
    .B2(_2086_),
    .X(_1139_));
 sky130_fd_sc_hd__or2_1 _4449_ (.A(net2057),
    .B(_2013_),
    .X(_2087_));
 sky130_fd_sc_hd__nor2_1 _4450_ (.A(_2014_),
    .B(net293),
    .Y(_2088_));
 sky130_fd_sc_hd__a22o_1 _4451_ (.A1(net2052),
    .A2(net293),
    .B1(_2087_),
    .B2(_2088_),
    .X(_1138_));
 sky130_fd_sc_hd__or2_1 _4452_ (.A(_1996_),
    .B(_2004_),
    .X(_2089_));
 sky130_fd_sc_hd__nor2_1 _4453_ (.A(net2057),
    .B(net293),
    .Y(_2090_));
 sky130_fd_sc_hd__a22o_1 _4454_ (.A1(net2055),
    .A2(net293),
    .B1(_2089_),
    .B2(_2090_),
    .X(_1137_));
 sky130_fd_sc_hd__or2_1 _4455_ (.A(_1987_),
    .B(_1995_),
    .X(_2091_));
 sky130_fd_sc_hd__nor2_1 _4456_ (.A(_1996_),
    .B(net294),
    .Y(_2092_));
 sky130_fd_sc_hd__a22o_1 _4457_ (.A1(net2059),
    .A2(net294),
    .B1(_2091_),
    .B2(_2092_),
    .X(_1136_));
 sky130_fd_sc_hd__a31o_1 _4458_ (.A1(_1960_),
    .A2(_1968_),
    .A3(_1978_),
    .B1(_1986_),
    .X(_2093_));
 sky130_fd_sc_hd__nor2_1 _4459_ (.A(_1987_),
    .B(net294),
    .Y(_2094_));
 sky130_fd_sc_hd__a22o_1 _4460_ (.A1(net2021),
    .A2(net294),
    .B1(_2093_),
    .B2(_2094_),
    .X(_1135_));
 sky130_fd_sc_hd__or2_1 _4461_ (.A(_1969_),
    .B(_1978_),
    .X(_2095_));
 sky130_fd_sc_hd__a21oi_1 _4462_ (.A1(_1969_),
    .A2(_1978_),
    .B1(net294),
    .Y(_2096_));
 sky130_fd_sc_hd__a22o_1 _4463_ (.A1(net1988),
    .A2(net294),
    .B1(_2095_),
    .B2(_2096_),
    .X(_1134_));
 sky130_fd_sc_hd__or2_1 _4464_ (.A(net2026),
    .B(_1968_),
    .X(_2097_));
 sky130_fd_sc_hd__nor2_1 _4465_ (.A(_1969_),
    .B(net295),
    .Y(_2098_));
 sky130_fd_sc_hd__a22o_1 _4466_ (.A1(net1874),
    .A2(net295),
    .B1(_2097_),
    .B2(_2098_),
    .X(_1133_));
 sky130_fd_sc_hd__a31o_1 _4467_ (.A1(_1932_),
    .A2(_1940_),
    .A3(_1949_),
    .B1(_1959_),
    .X(_2099_));
 sky130_fd_sc_hd__nor2_1 _4468_ (.A(_1960_),
    .B(net296),
    .Y(_2100_));
 sky130_fd_sc_hd__a22o_1 _4469_ (.A1(net2064),
    .A2(net296),
    .B1(_2099_),
    .B2(_2100_),
    .X(_1132_));
 sky130_fd_sc_hd__and2_1 _4470_ (.A(net2024),
    .B(net299),
    .X(_2101_));
 sky130_fd_sc_hd__or2_1 _4471_ (.A(_1941_),
    .B(_1949_),
    .X(_2102_));
 sky130_fd_sc_hd__a31o_1 _4472_ (.A1(_1950_),
    .A2(net284),
    .A3(_2102_),
    .B1(_2101_),
    .X(_1131_));
 sky130_fd_sc_hd__or2_1 _4473_ (.A(_1932_),
    .B(_1940_),
    .X(_2103_));
 sky130_fd_sc_hd__nor2_1 _4474_ (.A(_1941_),
    .B(net299),
    .Y(_2104_));
 sky130_fd_sc_hd__a22o_1 _4475_ (.A1(net2070),
    .A2(net299),
    .B1(_2103_),
    .B2(_2104_),
    .X(_1130_));
 sky130_fd_sc_hd__a21oi_1 _4476_ (.A1(_1914_),
    .A2(_1922_),
    .B1(_1931_),
    .Y(_2105_));
 sky130_fd_sc_hd__nor2_1 _4477_ (.A(_1932_),
    .B(_2105_),
    .Y(_2106_));
 sky130_fd_sc_hd__mux2_1 _4478_ (.A0(net2068),
    .A1(_2106_),
    .S(net285),
    .X(_1129_));
 sky130_fd_sc_hd__xor2_1 _4479_ (.A(_1914_),
    .B(_1922_),
    .X(_2107_));
 sky130_fd_sc_hd__mux2_1 _4480_ (.A0(net2023),
    .A1(_2107_),
    .S(net284),
    .X(_1128_));
 sky130_fd_sc_hd__or2_1 _4481_ (.A(_1905_),
    .B(_1913_),
    .X(_2108_));
 sky130_fd_sc_hd__nor2_1 _4482_ (.A(_1914_),
    .B(net297),
    .Y(_2109_));
 sky130_fd_sc_hd__a22o_1 _4483_ (.A1(net2015),
    .A2(net297),
    .B1(_2108_),
    .B2(_2109_),
    .X(_1127_));
 sky130_fd_sc_hd__nand2b_1 _4484_ (.A_N(_1904_),
    .B(net2028),
    .Y(_2110_));
 sky130_fd_sc_hd__nor2_1 _4485_ (.A(_1905_),
    .B(net297),
    .Y(_2111_));
 sky130_fd_sc_hd__a22o_1 _4486_ (.A1(net1989),
    .A2(net297),
    .B1(_2110_),
    .B2(_2111_),
    .X(_1126_));
 sky130_fd_sc_hd__and2_1 _4487_ (.A(net1971),
    .B(net297),
    .X(_2112_));
 sky130_fd_sc_hd__a31o_1 _4488_ (.A1(_1869_),
    .A2(_1877_),
    .A3(_1886_),
    .B1(_1894_),
    .X(_2113_));
 sky130_fd_sc_hd__a31o_1 _4489_ (.A1(net2028),
    .A2(net280),
    .A3(_2113_),
    .B1(_2112_),
    .X(_1125_));
 sky130_fd_sc_hd__xnor2_1 _4490_ (.A(_1878_),
    .B(_1886_),
    .Y(_2114_));
 sky130_fd_sc_hd__mux2_1 _4491_ (.A0(net2027),
    .A1(_2114_),
    .S(net282),
    .X(_1124_));
 sky130_fd_sc_hd__and2_1 _4492_ (.A(net2060),
    .B(net298),
    .X(_2115_));
 sky130_fd_sc_hd__or2_1 _4493_ (.A(_1869_),
    .B(_1877_),
    .X(_2116_));
 sky130_fd_sc_hd__a31o_1 _4494_ (.A1(_1878_),
    .A2(net280),
    .A3(_2116_),
    .B1(_2115_),
    .X(_1123_));
 sky130_fd_sc_hd__or2_1 _4495_ (.A(_1860_),
    .B(_1868_),
    .X(_2117_));
 sky130_fd_sc_hd__nor2_1 _4496_ (.A(_1869_),
    .B(net297),
    .Y(_2118_));
 sky130_fd_sc_hd__a22o_1 _4497_ (.A1(net2044),
    .A2(net297),
    .B1(_2117_),
    .B2(_2118_),
    .X(_1122_));
 sky130_fd_sc_hd__xnor2_1 _4498_ (.A(_1851_),
    .B(_1859_),
    .Y(_2119_));
 sky130_fd_sc_hd__mux2_1 _4499_ (.A0(net2013),
    .A1(_2119_),
    .S(net288),
    .X(_1121_));
 sky130_fd_sc_hd__and2_1 _4500_ (.A(net2061),
    .B(net300),
    .X(_2120_));
 sky130_fd_sc_hd__nand2b_1 _4501_ (.A_N(_1850_),
    .B(_1841_),
    .Y(_2121_));
 sky130_fd_sc_hd__a31o_1 _4502_ (.A1(_1851_),
    .A2(net287),
    .A3(_2121_),
    .B1(_2120_),
    .X(_1120_));
 sky130_fd_sc_hd__and2_1 _4503_ (.A(net2017),
    .B(net298),
    .X(_2122_));
 sky130_fd_sc_hd__nand2b_1 _4504_ (.A_N(_1840_),
    .B(_1832_),
    .Y(_2123_));
 sky130_fd_sc_hd__a31o_1 _4505_ (.A1(_1841_),
    .A2(net281),
    .A3(_2123_),
    .B1(_2122_),
    .X(_1119_));
 sky130_fd_sc_hd__and2_1 _4506_ (.A(net1992),
    .B(net299),
    .X(_2124_));
 sky130_fd_sc_hd__o21ai_1 _4507_ (.A1(_1813_),
    .A2(_1822_),
    .B1(_1831_),
    .Y(_2125_));
 sky130_fd_sc_hd__a31o_1 _4508_ (.A1(_1832_),
    .A2(net281),
    .A3(_2125_),
    .B1(_2124_),
    .X(_1118_));
 sky130_fd_sc_hd__xnor2_1 _4509_ (.A(_1813_),
    .B(_1821_),
    .Y(_2126_));
 sky130_fd_sc_hd__mux2_1 _4510_ (.A0(net1993),
    .A1(_2126_),
    .S(net281),
    .X(_1117_));
 sky130_fd_sc_hd__and2_1 _4511_ (.A(net2054),
    .B(net298),
    .X(_2127_));
 sky130_fd_sc_hd__a21o_1 _4512_ (.A1(_1799_),
    .A2(_1802_),
    .B1(_1812_),
    .X(_2128_));
 sky130_fd_sc_hd__a31o_1 _4513_ (.A1(_1813_),
    .A2(net281),
    .A3(_2128_),
    .B1(_2127_),
    .X(_1116_));
 sky130_fd_sc_hd__and2_1 _4514_ (.A(net2004),
    .B(net299),
    .X(_2129_));
 sky130_fd_sc_hd__or2_1 _4515_ (.A(_1799_),
    .B(_1802_),
    .X(_2130_));
 sky130_fd_sc_hd__a31o_1 _4516_ (.A1(_1804_),
    .A2(net281),
    .A3(_2130_),
    .B1(_2129_),
    .X(_1115_));
 sky130_fd_sc_hd__mux2_1 _4517_ (.A0(net2100),
    .A1(_1803_),
    .S(net276),
    .X(_1114_));
 sky130_fd_sc_hd__mux2_1 _4518_ (.A0(net2106),
    .A1(_2053_),
    .S(net272),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _4519_ (.A0(net2012),
    .A1(_2047_),
    .S(net271),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _4520_ (.A0(net1960),
    .A1(net2032),
    .S(net276),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _4521_ (.A0(net1850),
    .A1(_2031_),
    .S(net271),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _4522_ (.A0(net2179),
    .A1(_2022_),
    .S(net272),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _4523_ (.A0(net1713),
    .A1(net2053),
    .S(net274),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _4524_ (.A0(net796),
    .A1(net2056),
    .S(net272),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _4525_ (.A0(net1997),
    .A1(_1995_),
    .S(net274),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _4526_ (.A0(net929),
    .A1(_1986_),
    .S(net272),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _4527_ (.A0(net2119),
    .A1(_1978_),
    .S(net275),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _4528_ (.A0(net2095),
    .A1(_1968_),
    .S(net275),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _4529_ (.A0(net779),
    .A1(_1959_),
    .S(net271),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _4530_ (.A0(net1797),
    .A1(net2025),
    .S(net284),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _4531_ (.A0(net1943),
    .A1(_1940_),
    .S(net287),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _4532_ (.A0(net1944),
    .A1(net2079),
    .S(net285),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _4533_ (.A0(net2123),
    .A1(_1922_),
    .S(net280),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _4534_ (.A0(net1901),
    .A1(_1913_),
    .S(net287),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _4535_ (.A0(net2046),
    .A1(_1904_),
    .S(net279),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _4536_ (.A0(net809),
    .A1(_1894_),
    .S(net280),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _4537_ (.A0(net1780),
    .A1(_1886_),
    .S(net289),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _4538_ (.A0(net2011),
    .A1(_1877_),
    .S(net280),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _4539_ (.A0(net2088),
    .A1(_1868_),
    .S(net279),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _4540_ (.A0(net2069),
    .A1(_1859_),
    .S(net287),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _4541_ (.A0(net2242),
    .A1(_1850_),
    .S(net287),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _4542_ (.A0(net1417),
    .A1(_1840_),
    .S(net281),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _4543_ (.A0(net2035),
    .A1(_1830_),
    .S(net282),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _4544_ (.A0(net2117),
    .A1(_1821_),
    .S(net282),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _4545_ (.A0(net2120),
    .A1(_1812_),
    .S(net281),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _4546_ (.A0(net1995),
    .A1(_1799_),
    .S(net282),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _4547_ (.A0(net745),
    .A1(_1802_),
    .S(net276),
    .X(_0195_));
 sky130_fd_sc_hd__nand2b_2 _4548_ (.A_N(net2071),
    .B(net2144),
    .Y(_2131_));
 sky130_fd_sc_hd__nor3_1 _4549_ (.A(_1277_),
    .B(_1278_),
    .C(_2131_),
    .Y(_2132_));
 sky130_fd_sc_hd__or3_2 _4550_ (.A(_1277_),
    .B(_1278_),
    .C(_2131_),
    .X(_2133_));
 sky130_fd_sc_hd__and4bb_4 _4551_ (.A_N(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .B_N(net2048),
    .C(net2000),
    .D(net2071),
    .X(_2134_));
 sky130_fd_sc_hd__or4b_4 _4552_ (.A(net2124),
    .B(net2048),
    .C(_1278_),
    .D_N(net2071),
    .X(_2135_));
 sky130_fd_sc_hd__o21a_1 _4553_ (.A1(net2144),
    .A2(_2135_),
    .B1(_2133_),
    .X(_2136_));
 sky130_fd_sc_hd__or2_4 _4554_ (.A(net2048),
    .B(net2000),
    .X(_2137_));
 sky130_fd_sc_hd__o31a_1 _4555_ (.A1(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .A2(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .A3(_2137_),
    .B1(_2136_),
    .X(_3623_));
 sky130_fd_sc_hd__mux4_1 _4556_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ),
    .S0(net404),
    .S1(net394),
    .X(_2138_));
 sky130_fd_sc_hd__mux4_1 _4557_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ),
    .S0(net401),
    .S1(net394),
    .X(_2139_));
 sky130_fd_sc_hd__mux2_1 _4558_ (.A0(_2138_),
    .A1(_2139_),
    .S(net385),
    .X(_2140_));
 sky130_fd_sc_hd__mux4_1 _4559_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ),
    .S0(net401),
    .S1(net394),
    .X(_2141_));
 sky130_fd_sc_hd__mux4_1 _4560_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ),
    .S0(net404),
    .S1(net394),
    .X(_2142_));
 sky130_fd_sc_hd__mux2_1 _4561_ (.A0(_2142_),
    .A1(_2141_),
    .S(net385),
    .X(_2143_));
 sky130_fd_sc_hd__mux2_1 _4562_ (.A0(_2143_),
    .A1(_2140_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .X(_0000_));
 sky130_fd_sc_hd__mux4_1 _4563_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ),
    .S0(net404),
    .S1(net394),
    .X(_2144_));
 sky130_fd_sc_hd__mux4_1 _4564_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ),
    .S0(net404),
    .S1(net394),
    .X(_2145_));
 sky130_fd_sc_hd__mux2_1 _4565_ (.A0(_2144_),
    .A1(_2145_),
    .S(net385),
    .X(_2146_));
 sky130_fd_sc_hd__mux4_1 _4566_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ),
    .S0(net404),
    .S1(net394),
    .X(_2147_));
 sky130_fd_sc_hd__mux4_1 _4567_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ),
    .S0(net405),
    .S1(net395),
    .X(_2148_));
 sky130_fd_sc_hd__mux2_1 _4568_ (.A0(_2148_),
    .A1(_2147_),
    .S(net384),
    .X(_2149_));
 sky130_fd_sc_hd__mux2_1 _4569_ (.A0(_2149_),
    .A1(_2146_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .X(_0011_));
 sky130_fd_sc_hd__mux4_1 _4570_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ),
    .S0(net406),
    .S1(net391),
    .X(_2150_));
 sky130_fd_sc_hd__mux4_1 _4571_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ),
    .S0(net401),
    .S1(net391),
    .X(_2151_));
 sky130_fd_sc_hd__mux2_1 _4572_ (.A0(_2150_),
    .A1(_2151_),
    .S(net383),
    .X(_2152_));
 sky130_fd_sc_hd__mux4_1 _4573_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ),
    .S0(net406),
    .S1(net391),
    .X(_2153_));
 sky130_fd_sc_hd__mux4_1 _4574_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ),
    .S0(net406),
    .S1(net391),
    .X(_2154_));
 sky130_fd_sc_hd__mux2_1 _4575_ (.A0(_2154_),
    .A1(_2153_),
    .S(net383),
    .X(_2155_));
 sky130_fd_sc_hd__mux2_1 _4576_ (.A0(_2155_),
    .A1(_2152_),
    .S(net379),
    .X(_0022_));
 sky130_fd_sc_hd__mux4_1 _4577_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ),
    .S0(net404),
    .S1(net394),
    .X(_2156_));
 sky130_fd_sc_hd__mux4_1 _4578_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ),
    .S0(net404),
    .S1(net394),
    .X(_2157_));
 sky130_fd_sc_hd__mux2_1 _4579_ (.A0(_2156_),
    .A1(_2157_),
    .S(net385),
    .X(_2158_));
 sky130_fd_sc_hd__mux4_1 _4580_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ),
    .S0(net405),
    .S1(net394),
    .X(_2159_));
 sky130_fd_sc_hd__mux4_1 _4581_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ),
    .S0(net405),
    .S1(net395),
    .X(_2160_));
 sky130_fd_sc_hd__mux2_1 _4582_ (.A0(_2160_),
    .A1(_2159_),
    .S(net385),
    .X(_2161_));
 sky130_fd_sc_hd__mux2_1 _4583_ (.A0(_2161_),
    .A1(_2158_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .X(_0025_));
 sky130_fd_sc_hd__mux4_1 _4584_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ),
    .S0(net403),
    .S1(net393),
    .X(_2162_));
 sky130_fd_sc_hd__mux4_1 _4585_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ),
    .S0(net403),
    .S1(net393),
    .X(_2163_));
 sky130_fd_sc_hd__mux2_1 _4586_ (.A0(_2162_),
    .A1(_2163_),
    .S(net384),
    .X(_2164_));
 sky130_fd_sc_hd__mux4_1 _4587_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ),
    .S0(net403),
    .S1(net393),
    .X(_2165_));
 sky130_fd_sc_hd__mux4_1 _4588_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ),
    .S0(net406),
    .S1(net393),
    .X(_2166_));
 sky130_fd_sc_hd__mux2_1 _4589_ (.A0(_2166_),
    .A1(_2165_),
    .S(net384),
    .X(_2167_));
 sky130_fd_sc_hd__mux2_1 _4590_ (.A0(_2167_),
    .A1(_2164_),
    .S(net379),
    .X(_0026_));
 sky130_fd_sc_hd__mux4_1 _4591_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ),
    .S0(net402),
    .S1(net391),
    .X(_2168_));
 sky130_fd_sc_hd__mux4_1 _4592_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ),
    .S0(net403),
    .S1(net392),
    .X(_2169_));
 sky130_fd_sc_hd__mux2_1 _4593_ (.A0(_2168_),
    .A1(_2169_),
    .S(net384),
    .X(_2170_));
 sky130_fd_sc_hd__mux4_1 _4594_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ),
    .S0(net403),
    .S1(net392),
    .X(_2171_));
 sky130_fd_sc_hd__mux4_1 _4595_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ),
    .S0(net403),
    .S1(net392),
    .X(_2172_));
 sky130_fd_sc_hd__mux2_1 _4596_ (.A0(_2172_),
    .A1(_2171_),
    .S(net384),
    .X(_2173_));
 sky130_fd_sc_hd__mux2_1 _4597_ (.A0(_2173_),
    .A1(_2170_),
    .S(net379),
    .X(_0027_));
 sky130_fd_sc_hd__mux4_1 _4598_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ),
    .S0(net401),
    .S1(net391),
    .X(_2174_));
 sky130_fd_sc_hd__mux4_1 _4599_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ),
    .S0(net401),
    .S1(net391),
    .X(_2175_));
 sky130_fd_sc_hd__mux2_1 _4600_ (.A0(_2174_),
    .A1(_2175_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ),
    .X(_2176_));
 sky130_fd_sc_hd__mux4_1 _4601_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ),
    .S0(net401),
    .S1(net391),
    .X(_2177_));
 sky130_fd_sc_hd__mux4_1 _4602_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ),
    .S0(net401),
    .S1(net391),
    .X(_2178_));
 sky130_fd_sc_hd__mux2_1 _4603_ (.A0(_2178_),
    .A1(_2177_),
    .S(net383),
    .X(_2179_));
 sky130_fd_sc_hd__mux2_1 _4604_ (.A0(_2179_),
    .A1(_2176_),
    .S(net379),
    .X(_0028_));
 sky130_fd_sc_hd__mux4_1 _4605_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ),
    .S0(net402),
    .S1(net390),
    .X(_2180_));
 sky130_fd_sc_hd__mux4_1 _4606_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ),
    .S0(net402),
    .S1(net390),
    .X(_2181_));
 sky130_fd_sc_hd__mux2_1 _4607_ (.A0(_2180_),
    .A1(_2181_),
    .S(net383),
    .X(_2182_));
 sky130_fd_sc_hd__mux4_1 _4608_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ),
    .S0(net401),
    .S1(net390),
    .X(_2183_));
 sky130_fd_sc_hd__mux4_1 _4609_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ),
    .S0(net401),
    .S1(net390),
    .X(_2184_));
 sky130_fd_sc_hd__mux2_1 _4610_ (.A0(_2184_),
    .A1(_2183_),
    .S(net383),
    .X(_2185_));
 sky130_fd_sc_hd__mux2_1 _4611_ (.A0(_2185_),
    .A1(_2182_),
    .S(net379),
    .X(_0029_));
 sky130_fd_sc_hd__mux4_1 _4612_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ),
    .S0(net402),
    .S1(net390),
    .X(_2186_));
 sky130_fd_sc_hd__mux4_1 _4613_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ),
    .S0(net402),
    .S1(net390),
    .X(_2187_));
 sky130_fd_sc_hd__mux2_1 _4614_ (.A0(_2186_),
    .A1(_2187_),
    .S(net383),
    .X(_2188_));
 sky130_fd_sc_hd__mux4_1 _4615_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ),
    .S0(net402),
    .S1(net390),
    .X(_2189_));
 sky130_fd_sc_hd__mux4_1 _4616_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ),
    .S0(net402),
    .S1(net391),
    .X(_2190_));
 sky130_fd_sc_hd__mux2_1 _4617_ (.A0(_2190_),
    .A1(_2189_),
    .S(net383),
    .X(_2191_));
 sky130_fd_sc_hd__mux2_1 _4618_ (.A0(_2191_),
    .A1(_2188_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .X(_0030_));
 sky130_fd_sc_hd__mux4_1 _4619_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ),
    .S0(net405),
    .S1(net395),
    .X(_2192_));
 sky130_fd_sc_hd__mux4_1 _4620_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ),
    .S0(net405),
    .S1(net394),
    .X(_2193_));
 sky130_fd_sc_hd__mux2_1 _4621_ (.A0(_2192_),
    .A1(_2193_),
    .S(net385),
    .X(_2194_));
 sky130_fd_sc_hd__mux4_1 _4622_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ),
    .S0(net405),
    .S1(net394),
    .X(_2195_));
 sky130_fd_sc_hd__mux4_1 _4623_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ),
    .S0(net405),
    .S1(net394),
    .X(_2196_));
 sky130_fd_sc_hd__mux2_1 _4624_ (.A0(_2196_),
    .A1(_2195_),
    .S(net385),
    .X(_2197_));
 sky130_fd_sc_hd__mux2_1 _4625_ (.A0(_2197_),
    .A1(_2194_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .X(_0031_));
 sky130_fd_sc_hd__mux4_1 _4626_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ),
    .S0(net403),
    .S1(net392),
    .X(_2198_));
 sky130_fd_sc_hd__mux4_1 _4627_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ),
    .S0(net403),
    .S1(net392),
    .X(_2199_));
 sky130_fd_sc_hd__mux2_1 _4628_ (.A0(_2198_),
    .A1(_2199_),
    .S(net384),
    .X(_2200_));
 sky130_fd_sc_hd__mux4_1 _4629_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ),
    .S0(net402),
    .S1(net390),
    .X(_2201_));
 sky130_fd_sc_hd__mux4_1 _4630_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ),
    .S0(net402),
    .S1(net390),
    .X(_2202_));
 sky130_fd_sc_hd__mux2_1 _4631_ (.A0(_2202_),
    .A1(_2201_),
    .S(net383),
    .X(_2203_));
 sky130_fd_sc_hd__mux2_1 _4632_ (.A0(_2203_),
    .A1(_2200_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .X(_0001_));
 sky130_fd_sc_hd__mux4_1 _4633_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ),
    .S0(net397),
    .S1(net387),
    .X(_2204_));
 sky130_fd_sc_hd__mux4_1 _4634_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ),
    .S0(net399),
    .S1(net388),
    .X(_2205_));
 sky130_fd_sc_hd__mux2_1 _4635_ (.A0(_2204_),
    .A1(_2205_),
    .S(net382),
    .X(_2206_));
 sky130_fd_sc_hd__mux4_1 _4636_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ),
    .S0(net399),
    .S1(net388),
    .X(_2207_));
 sky130_fd_sc_hd__mux4_1 _4637_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ),
    .S0(net399),
    .S1(net388),
    .X(_2208_));
 sky130_fd_sc_hd__mux2_1 _4638_ (.A0(_2208_),
    .A1(_2207_),
    .S(net382),
    .X(_2209_));
 sky130_fd_sc_hd__mux2_1 _4639_ (.A0(_2209_),
    .A1(_2206_),
    .S(net380),
    .X(_0002_));
 sky130_fd_sc_hd__mux4_1 _4640_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ),
    .S0(net403),
    .S1(net392),
    .X(_2210_));
 sky130_fd_sc_hd__mux4_1 _4641_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ),
    .S0(net406),
    .S1(net392),
    .X(_2211_));
 sky130_fd_sc_hd__mux2_1 _4642_ (.A0(_2210_),
    .A1(_2211_),
    .S(net384),
    .X(_2212_));
 sky130_fd_sc_hd__mux4_1 _4643_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ),
    .S0(net403),
    .S1(net393),
    .X(_2213_));
 sky130_fd_sc_hd__mux4_1 _4644_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ),
    .S0(net406),
    .S1(net393),
    .X(_2214_));
 sky130_fd_sc_hd__mux2_1 _4645_ (.A0(_2214_),
    .A1(_2213_),
    .S(net384),
    .X(_2215_));
 sky130_fd_sc_hd__mux2_1 _4646_ (.A0(_2215_),
    .A1(_2212_),
    .S(net379),
    .X(_0003_));
 sky130_fd_sc_hd__mux4_1 _4647_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ),
    .S0(net399),
    .S1(net389),
    .X(_2216_));
 sky130_fd_sc_hd__mux4_1 _4648_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ),
    .S0(net399),
    .S1(net388),
    .X(_2217_));
 sky130_fd_sc_hd__mux2_1 _4649_ (.A0(_2216_),
    .A1(_2217_),
    .S(net382),
    .X(_2218_));
 sky130_fd_sc_hd__mux4_1 _4650_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ),
    .S0(net399),
    .S1(net388),
    .X(_2219_));
 sky130_fd_sc_hd__mux4_1 _4651_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ),
    .S0(net399),
    .S1(net388),
    .X(_2220_));
 sky130_fd_sc_hd__mux2_1 _4652_ (.A0(_2220_),
    .A1(_2219_),
    .S(net382),
    .X(_2221_));
 sky130_fd_sc_hd__mux2_1 _4653_ (.A0(_2221_),
    .A1(_2218_),
    .S(net380),
    .X(_0004_));
 sky130_fd_sc_hd__mux4_1 _4654_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ),
    .S0(net402),
    .S1(net390),
    .X(_2222_));
 sky130_fd_sc_hd__mux4_1 _4655_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ),
    .S0(net402),
    .S1(net390),
    .X(_2223_));
 sky130_fd_sc_hd__mux2_1 _4656_ (.A0(_2222_),
    .A1(_2223_),
    .S(net383),
    .X(_2224_));
 sky130_fd_sc_hd__mux4_1 _4657_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ),
    .S0(net402),
    .S1(net390),
    .X(_2225_));
 sky130_fd_sc_hd__mux4_1 _4658_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ),
    .S0(net402),
    .S1(net390),
    .X(_2226_));
 sky130_fd_sc_hd__mux2_1 _4659_ (.A0(_2226_),
    .A1(_2225_),
    .S(net383),
    .X(_2227_));
 sky130_fd_sc_hd__mux2_1 _4660_ (.A0(_2227_),
    .A1(_2224_),
    .S(net379),
    .X(_0005_));
 sky130_fd_sc_hd__mux4_1 _4661_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ),
    .S0(net403),
    .S1(net392),
    .X(_2228_));
 sky130_fd_sc_hd__mux4_1 _4662_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ),
    .S0(net403),
    .S1(net392),
    .X(_2229_));
 sky130_fd_sc_hd__mux2_1 _4663_ (.A0(_2228_),
    .A1(_2229_),
    .S(net384),
    .X(_2230_));
 sky130_fd_sc_hd__mux4_1 _4664_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ),
    .S0(net403),
    .S1(net392),
    .X(_2231_));
 sky130_fd_sc_hd__mux4_1 _4665_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ),
    .S0(net403),
    .S1(net392),
    .X(_2232_));
 sky130_fd_sc_hd__mux2_1 _4666_ (.A0(_2232_),
    .A1(_2231_),
    .S(net384),
    .X(_2233_));
 sky130_fd_sc_hd__mux2_1 _4667_ (.A0(_2233_),
    .A1(_2230_),
    .S(net379),
    .X(_0006_));
 sky130_fd_sc_hd__mux4_1 _4668_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ),
    .S0(net399),
    .S1(net389),
    .X(_2234_));
 sky130_fd_sc_hd__mux4_1 _4669_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ),
    .S0(net399),
    .S1(net389),
    .X(_2235_));
 sky130_fd_sc_hd__mux2_1 _4670_ (.A0(_2234_),
    .A1(_2235_),
    .S(net382),
    .X(_2236_));
 sky130_fd_sc_hd__mux4_1 _4671_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ),
    .S0(net399),
    .S1(net388),
    .X(_2237_));
 sky130_fd_sc_hd__mux4_1 _4672_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ),
    .S0(net400),
    .S1(net388),
    .X(_2238_));
 sky130_fd_sc_hd__mux2_1 _4673_ (.A0(_2238_),
    .A1(_2237_),
    .S(net382),
    .X(_2239_));
 sky130_fd_sc_hd__mux2_1 _4674_ (.A0(_2239_),
    .A1(_2236_),
    .S(net380),
    .X(_0007_));
 sky130_fd_sc_hd__mux4_1 _4675_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ),
    .S0(net398),
    .S1(net387),
    .X(_2240_));
 sky130_fd_sc_hd__mux4_1 _4676_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ),
    .S0(net398),
    .S1(net387),
    .X(_2241_));
 sky130_fd_sc_hd__mux2_1 _4677_ (.A0(_2240_),
    .A1(_2241_),
    .S(net381),
    .X(_2242_));
 sky130_fd_sc_hd__mux4_1 _4678_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ),
    .S0(net398),
    .S1(net387),
    .X(_2243_));
 sky130_fd_sc_hd__mux4_1 _4679_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ),
    .S0(net398),
    .S1(net387),
    .X(_2244_));
 sky130_fd_sc_hd__mux2_1 _4680_ (.A0(_2244_),
    .A1(_2243_),
    .S(net381),
    .X(_2245_));
 sky130_fd_sc_hd__mux2_1 _4681_ (.A0(_2245_),
    .A1(_2242_),
    .S(net380),
    .X(_0008_));
 sky130_fd_sc_hd__mux4_1 _4682_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ),
    .S0(net404),
    .S1(net392),
    .X(_2246_));
 sky130_fd_sc_hd__mux4_1 _4683_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ),
    .S0(net404),
    .S1(net392),
    .X(_2247_));
 sky130_fd_sc_hd__mux2_1 _4684_ (.A0(_2246_),
    .A1(_2247_),
    .S(net384),
    .X(_2248_));
 sky130_fd_sc_hd__mux4_1 _4685_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ),
    .S0(net404),
    .S1(net394),
    .X(_2249_));
 sky130_fd_sc_hd__mux4_1 _4686_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ),
    .S0(net404),
    .S1(net394),
    .X(_2250_));
 sky130_fd_sc_hd__mux2_1 _4687_ (.A0(_2250_),
    .A1(_2249_),
    .S(net385),
    .X(_2251_));
 sky130_fd_sc_hd__mux2_1 _4688_ (.A0(_2251_),
    .A1(_2248_),
    .S(net379),
    .X(_0009_));
 sky130_fd_sc_hd__mux4_1 _4689_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ),
    .S0(net400),
    .S1(net389),
    .X(_2252_));
 sky130_fd_sc_hd__mux4_1 _4690_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ),
    .S0(net400),
    .S1(net389),
    .X(_2253_));
 sky130_fd_sc_hd__mux2_1 _4691_ (.A0(_2252_),
    .A1(_2253_),
    .S(net382),
    .X(_2254_));
 sky130_fd_sc_hd__mux4_1 _4692_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ),
    .S0(net400),
    .S1(net389),
    .X(_2255_));
 sky130_fd_sc_hd__mux4_1 _4693_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ),
    .S0(net400),
    .S1(net389),
    .X(_2256_));
 sky130_fd_sc_hd__mux2_1 _4694_ (.A0(_2256_),
    .A1(_2255_),
    .S(net382),
    .X(_2257_));
 sky130_fd_sc_hd__mux2_1 _4695_ (.A0(_2257_),
    .A1(_2254_),
    .S(net380),
    .X(_0010_));
 sky130_fd_sc_hd__mux4_1 _4696_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ),
    .S0(net396),
    .S1(net386),
    .X(_2258_));
 sky130_fd_sc_hd__mux4_1 _4697_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ),
    .S0(net397),
    .S1(net386),
    .X(_2259_));
 sky130_fd_sc_hd__mux2_1 _4698_ (.A0(_2258_),
    .A1(_2259_),
    .S(net381),
    .X(_2260_));
 sky130_fd_sc_hd__mux4_1 _4699_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ),
    .S0(net396),
    .S1(net386),
    .X(_2261_));
 sky130_fd_sc_hd__mux4_1 _4700_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ),
    .S0(net396),
    .S1(net386),
    .X(_2262_));
 sky130_fd_sc_hd__mux2_1 _4701_ (.A0(_2262_),
    .A1(_2261_),
    .S(net381),
    .X(_2263_));
 sky130_fd_sc_hd__mux2_1 _4702_ (.A0(_2263_),
    .A1(_2260_),
    .S(net380),
    .X(_0012_));
 sky130_fd_sc_hd__mux4_1 _4703_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ),
    .S0(net397),
    .S1(net388),
    .X(_2264_));
 sky130_fd_sc_hd__mux4_1 _4704_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ),
    .S0(net397),
    .S1(net388),
    .X(_2265_));
 sky130_fd_sc_hd__mux2_1 _4705_ (.A0(_2264_),
    .A1(_2265_),
    .S(net382),
    .X(_2266_));
 sky130_fd_sc_hd__mux4_1 _4706_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ),
    .S0(net397),
    .S1(net387),
    .X(_2267_));
 sky130_fd_sc_hd__mux4_1 _4707_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ),
    .S0(net397),
    .S1(net387),
    .X(_2268_));
 sky130_fd_sc_hd__mux2_1 _4708_ (.A0(_2268_),
    .A1(_2267_),
    .S(net381),
    .X(_2269_));
 sky130_fd_sc_hd__mux2_1 _4709_ (.A0(_2269_),
    .A1(_2266_),
    .S(net380),
    .X(_0013_));
 sky130_fd_sc_hd__mux4_1 _4710_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ),
    .S0(net401),
    .S1(net391),
    .X(_2270_));
 sky130_fd_sc_hd__mux4_1 _4711_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ),
    .S0(net401),
    .S1(net391),
    .X(_2271_));
 sky130_fd_sc_hd__mux2_1 _4712_ (.A0(_2270_),
    .A1(_2271_),
    .S(net383),
    .X(_2272_));
 sky130_fd_sc_hd__mux4_1 _4713_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ),
    .S0(net401),
    .S1(net391),
    .X(_2273_));
 sky130_fd_sc_hd__mux4_1 _4714_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ),
    .S0(net401),
    .S1(net391),
    .X(_2274_));
 sky130_fd_sc_hd__mux2_1 _4715_ (.A0(_2274_),
    .A1(_2273_),
    .S(net383),
    .X(_2275_));
 sky130_fd_sc_hd__mux2_1 _4716_ (.A0(_2275_),
    .A1(_2272_),
    .S(net379),
    .X(_0014_));
 sky130_fd_sc_hd__mux4_1 _4717_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ),
    .S0(net396),
    .S1(net387),
    .X(_2276_));
 sky130_fd_sc_hd__mux4_1 _4718_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ),
    .S0(net397),
    .S1(net386),
    .X(_2277_));
 sky130_fd_sc_hd__mux2_1 _4719_ (.A0(_2276_),
    .A1(_2277_),
    .S(net381),
    .X(_2278_));
 sky130_fd_sc_hd__mux4_1 _4720_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ),
    .S0(net396),
    .S1(net386),
    .X(_2279_));
 sky130_fd_sc_hd__mux4_1 _4721_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ),
    .S0(net396),
    .S1(net386),
    .X(_2280_));
 sky130_fd_sc_hd__mux2_1 _4722_ (.A0(_2280_),
    .A1(_2279_),
    .S(net381),
    .X(_2281_));
 sky130_fd_sc_hd__mux2_1 _4723_ (.A0(_2281_),
    .A1(_2278_),
    .S(net380),
    .X(_0015_));
 sky130_fd_sc_hd__mux4_1 _4724_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ),
    .S0(net404),
    .S1(net395),
    .X(_2282_));
 sky130_fd_sc_hd__mux4_1 _4725_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ),
    .S0(net405),
    .S1(net394),
    .X(_2283_));
 sky130_fd_sc_hd__mux2_1 _4726_ (.A0(_2282_),
    .A1(_2283_),
    .S(net384),
    .X(_2284_));
 sky130_fd_sc_hd__mux4_1 _4727_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ),
    .S0(net404),
    .S1(net392),
    .X(_2285_));
 sky130_fd_sc_hd__mux4_1 _4728_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ),
    .S0(net404),
    .S1(net395),
    .X(_2286_));
 sky130_fd_sc_hd__mux2_1 _4729_ (.A0(_2286_),
    .A1(_2285_),
    .S(net384),
    .X(_2287_));
 sky130_fd_sc_hd__mux2_1 _4730_ (.A0(_2287_),
    .A1(_2284_),
    .S(net379),
    .X(_0016_));
 sky130_fd_sc_hd__mux4_1 _4731_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ),
    .S0(net396),
    .S1(net387),
    .X(_2288_));
 sky130_fd_sc_hd__mux4_1 _4732_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ),
    .S0(net397),
    .S1(net386),
    .X(_2289_));
 sky130_fd_sc_hd__mux2_1 _4733_ (.A0(_2288_),
    .A1(_2289_),
    .S(net381),
    .X(_2290_));
 sky130_fd_sc_hd__mux4_1 _4734_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ),
    .S0(net396),
    .S1(net386),
    .X(_2291_));
 sky130_fd_sc_hd__mux4_1 _4735_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ),
    .S0(net396),
    .S1(net386),
    .X(_2292_));
 sky130_fd_sc_hd__mux2_1 _4736_ (.A0(_2292_),
    .A1(_2291_),
    .S(net381),
    .X(_2293_));
 sky130_fd_sc_hd__mux2_1 _4737_ (.A0(_2293_),
    .A1(_2290_),
    .S(net380),
    .X(_0017_));
 sky130_fd_sc_hd__mux4_1 _4738_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ),
    .S0(net397),
    .S1(net386),
    .X(_2294_));
 sky130_fd_sc_hd__mux4_1 _4739_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ),
    .S0(net397),
    .S1(net386),
    .X(_2295_));
 sky130_fd_sc_hd__mux2_1 _4740_ (.A0(_2294_),
    .A1(_2295_),
    .S(net381),
    .X(_2296_));
 sky130_fd_sc_hd__mux4_1 _4741_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ),
    .S0(net396),
    .S1(net386),
    .X(_2297_));
 sky130_fd_sc_hd__mux4_1 _4742_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ),
    .S0(net396),
    .S1(net386),
    .X(_2298_));
 sky130_fd_sc_hd__mux2_1 _4743_ (.A0(_2298_),
    .A1(_2297_),
    .S(net381),
    .X(_2299_));
 sky130_fd_sc_hd__mux2_1 _4744_ (.A0(_2299_),
    .A1(_2296_),
    .S(net380),
    .X(_0018_));
 sky130_fd_sc_hd__mux4_1 _4745_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ),
    .S0(net401),
    .S1(net391),
    .X(_2300_));
 sky130_fd_sc_hd__mux4_1 _4746_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ),
    .S0(net399),
    .S1(net389),
    .X(_2301_));
 sky130_fd_sc_hd__mux2_1 _4747_ (.A0(_2300_),
    .A1(_2301_),
    .S(net383),
    .X(_2302_));
 sky130_fd_sc_hd__mux4_1 _4748_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ),
    .S0(net401),
    .S1(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ),
    .X(_2303_));
 sky130_fd_sc_hd__mux4_1 _4749_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ),
    .S0(net399),
    .S1(net388),
    .X(_2304_));
 sky130_fd_sc_hd__mux2_1 _4750_ (.A0(_2304_),
    .A1(_2303_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ),
    .X(_2305_));
 sky130_fd_sc_hd__mux2_1 _4751_ (.A0(_2305_),
    .A1(_2302_),
    .S(net379),
    .X(_0019_));
 sky130_fd_sc_hd__mux4_1 _4752_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ),
    .S0(net396),
    .S1(net386),
    .X(_2306_));
 sky130_fd_sc_hd__mux4_1 _4753_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ),
    .S0(net397),
    .S1(net388),
    .X(_2307_));
 sky130_fd_sc_hd__mux2_1 _4754_ (.A0(_2306_),
    .A1(_2307_),
    .S(net381),
    .X(_2308_));
 sky130_fd_sc_hd__mux4_1 _4755_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ),
    .S0(net396),
    .S1(net389),
    .X(_2309_));
 sky130_fd_sc_hd__mux4_1 _4756_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ),
    .S0(net397),
    .S1(net387),
    .X(_2310_));
 sky130_fd_sc_hd__mux2_1 _4757_ (.A0(_2310_),
    .A1(_2309_),
    .S(net382),
    .X(_2311_));
 sky130_fd_sc_hd__mux2_1 _4758_ (.A0(_2311_),
    .A1(_2308_),
    .S(net380),
    .X(_0020_));
 sky130_fd_sc_hd__mux4_1 _4759_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ),
    .S0(net396),
    .S1(net387),
    .X(_2312_));
 sky130_fd_sc_hd__mux4_1 _4760_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ),
    .S0(net397),
    .S1(net387),
    .X(_2313_));
 sky130_fd_sc_hd__mux2_1 _4761_ (.A0(_2312_),
    .A1(_2313_),
    .S(net381),
    .X(_2314_));
 sky130_fd_sc_hd__mux4_1 _4762_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ),
    .S0(net396),
    .S1(net387),
    .X(_2315_));
 sky130_fd_sc_hd__mux4_1 _4763_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ),
    .S0(net396),
    .S1(net387),
    .X(_2316_));
 sky130_fd_sc_hd__mux2_1 _4764_ (.A0(_2316_),
    .A1(_2315_),
    .S(net381),
    .X(_2317_));
 sky130_fd_sc_hd__mux2_1 _4765_ (.A0(_2317_),
    .A1(_2314_),
    .S(net380),
    .X(_0021_));
 sky130_fd_sc_hd__mux4_1 _4766_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ),
    .S0(net404),
    .S1(net392),
    .X(_2318_));
 sky130_fd_sc_hd__mux4_1 _4767_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ),
    .S0(net404),
    .S1(net392),
    .X(_2319_));
 sky130_fd_sc_hd__mux2_1 _4768_ (.A0(_2318_),
    .A1(_2319_),
    .S(net384),
    .X(_2320_));
 sky130_fd_sc_hd__mux4_1 _4769_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ),
    .S0(net403),
    .S1(net393),
    .X(_2321_));
 sky130_fd_sc_hd__mux4_1 _4770_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ),
    .S0(net403),
    .S1(net393),
    .X(_2322_));
 sky130_fd_sc_hd__mux2_1 _4771_ (.A0(_2322_),
    .A1(_2321_),
    .S(net384),
    .X(_2323_));
 sky130_fd_sc_hd__mux2_1 _4772_ (.A0(_2323_),
    .A1(_2320_),
    .S(net379),
    .X(_0023_));
 sky130_fd_sc_hd__mux4_1 _4773_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ),
    .S0(net399),
    .S1(net388),
    .X(_2324_));
 sky130_fd_sc_hd__mux4_1 _4774_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ),
    .S0(net399),
    .S1(net388),
    .X(_2325_));
 sky130_fd_sc_hd__mux2_1 _4775_ (.A0(_2324_),
    .A1(_2325_),
    .S(net381),
    .X(_2326_));
 sky130_fd_sc_hd__mux4_1 _4776_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ),
    .S0(net399),
    .S1(net388),
    .X(_2327_));
 sky130_fd_sc_hd__mux4_1 _4777_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ),
    .S0(net399),
    .S1(net388),
    .X(_2328_));
 sky130_fd_sc_hd__mux2_1 _4778_ (.A0(_2328_),
    .A1(_2327_),
    .S(net382),
    .X(_2329_));
 sky130_fd_sc_hd__mux2_1 _4779_ (.A0(_2329_),
    .A1(_2326_),
    .S(net380),
    .X(_0024_));
 sky130_fd_sc_hd__mux4_1 _4780_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ),
    .S0(net433),
    .S1(net423),
    .X(_2330_));
 sky130_fd_sc_hd__mux4_1 _4781_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ),
    .S0(net430),
    .S1(net421),
    .X(_2331_));
 sky130_fd_sc_hd__mux2_1 _4782_ (.A0(_2330_),
    .A1(_2331_),
    .S(net412),
    .X(_2332_));
 sky130_fd_sc_hd__mux4_1 _4783_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ),
    .S0(net430),
    .S1(net421),
    .X(_2333_));
 sky130_fd_sc_hd__mux4_1 _4784_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ),
    .S0(net433),
    .S1(net423),
    .X(_2334_));
 sky130_fd_sc_hd__mux2_1 _4785_ (.A0(_2334_),
    .A1(_2333_),
    .S(net412),
    .X(_2335_));
 sky130_fd_sc_hd__mux2_1 _4786_ (.A0(_2335_),
    .A1(_2332_),
    .S(net407),
    .X(_0032_));
 sky130_fd_sc_hd__mux4_1 _4787_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ),
    .S0(net433),
    .S1(net423),
    .X(_2336_));
 sky130_fd_sc_hd__mux4_1 _4788_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ),
    .S0(net433),
    .S1(net423),
    .X(_2337_));
 sky130_fd_sc_hd__mux2_1 _4789_ (.A0(_2336_),
    .A1(_2337_),
    .S(net413),
    .X(_2338_));
 sky130_fd_sc_hd__mux4_1 _4790_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ),
    .S0(net433),
    .S1(net423),
    .X(_2339_));
 sky130_fd_sc_hd__mux4_1 _4791_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ),
    .S0(net434),
    .S1(net424),
    .X(_2340_));
 sky130_fd_sc_hd__mux2_1 _4792_ (.A0(_2340_),
    .A1(_2339_),
    .S(net413),
    .X(_2341_));
 sky130_fd_sc_hd__mux2_1 _4793_ (.A0(_2341_),
    .A1(_2338_),
    .S(net407),
    .X(_0043_));
 sky130_fd_sc_hd__mux4_1 _4794_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ),
    .S0(net430),
    .S1(net421),
    .X(_2342_));
 sky130_fd_sc_hd__mux4_1 _4795_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ),
    .S0(net430),
    .S1(net421),
    .X(_2343_));
 sky130_fd_sc_hd__mux2_1 _4796_ (.A0(_2342_),
    .A1(_2343_),
    .S(net412),
    .X(_2344_));
 sky130_fd_sc_hd__mux4_1 _4797_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ),
    .S0(net430),
    .S1(net421),
    .X(_2345_));
 sky130_fd_sc_hd__mux4_1 _4798_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ),
    .S0(net430),
    .S1(net421),
    .X(_2346_));
 sky130_fd_sc_hd__mux2_1 _4799_ (.A0(_2346_),
    .A1(_2345_),
    .S(net412),
    .X(_2347_));
 sky130_fd_sc_hd__mux2_1 _4800_ (.A0(_2347_),
    .A1(_2344_),
    .S(net407),
    .X(_0054_));
 sky130_fd_sc_hd__mux4_1 _4801_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ),
    .S0(net433),
    .S1(net423),
    .X(_2348_));
 sky130_fd_sc_hd__mux4_1 _4802_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ),
    .S0(net433),
    .S1(net423),
    .X(_2349_));
 sky130_fd_sc_hd__mux2_1 _4803_ (.A0(_2348_),
    .A1(_2349_),
    .S(net412),
    .X(_2350_));
 sky130_fd_sc_hd__mux4_1 _4804_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ),
    .S0(net434),
    .S1(net423),
    .X(_2351_));
 sky130_fd_sc_hd__mux4_1 _4805_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ),
    .S0(net433),
    .S1(net423),
    .X(_2352_));
 sky130_fd_sc_hd__mux2_1 _4806_ (.A0(_2352_),
    .A1(_2351_),
    .S(net413),
    .X(_2353_));
 sky130_fd_sc_hd__mux2_1 _4807_ (.A0(_2353_),
    .A1(_2350_),
    .S(net407),
    .X(_0057_));
 sky130_fd_sc_hd__mux4_1 _4808_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ),
    .S0(net432),
    .S1(net422),
    .X(_2354_));
 sky130_fd_sc_hd__mux4_1 _4809_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ),
    .S0(net432),
    .S1(net424),
    .X(_2355_));
 sky130_fd_sc_hd__mux2_1 _4810_ (.A0(_2354_),
    .A1(_2355_),
    .S(net413),
    .X(_2356_));
 sky130_fd_sc_hd__mux4_1 _4811_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ),
    .S0(net431),
    .S1(net424),
    .X(_2357_));
 sky130_fd_sc_hd__mux4_1 _4812_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ),
    .S0(net431),
    .S1(net422),
    .X(_2358_));
 sky130_fd_sc_hd__mux2_1 _4813_ (.A0(_2358_),
    .A1(_2357_),
    .S(net412),
    .X(_2359_));
 sky130_fd_sc_hd__mux2_1 _4814_ (.A0(_2359_),
    .A1(_2356_),
    .S(net407),
    .X(_0058_));
 sky130_fd_sc_hd__mux4_1 _4815_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ),
    .S0(net430),
    .S1(net421),
    .X(_2360_));
 sky130_fd_sc_hd__mux4_1 _4816_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ),
    .S0(net431),
    .S1(net422),
    .X(_2361_));
 sky130_fd_sc_hd__mux2_1 _4817_ (.A0(_2360_),
    .A1(_2361_),
    .S(net412),
    .X(_2362_));
 sky130_fd_sc_hd__mux4_1 _4818_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ),
    .S0(net431),
    .S1(net422),
    .X(_2363_));
 sky130_fd_sc_hd__mux4_1 _4819_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ),
    .S0(net431),
    .S1(net422),
    .X(_2364_));
 sky130_fd_sc_hd__mux2_1 _4820_ (.A0(_2364_),
    .A1(_2363_),
    .S(net412),
    .X(_2365_));
 sky130_fd_sc_hd__mux2_1 _4821_ (.A0(_2365_),
    .A1(_2362_),
    .S(net407),
    .X(_0059_));
 sky130_fd_sc_hd__mux4_1 _4822_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ),
    .S0(net430),
    .S1(net421),
    .X(_2366_));
 sky130_fd_sc_hd__mux4_1 _4823_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ),
    .S0(net430),
    .S1(net421),
    .X(_2367_));
 sky130_fd_sc_hd__mux2_1 _4824_ (.A0(_2366_),
    .A1(_2367_),
    .S(net411),
    .X(_2368_));
 sky130_fd_sc_hd__mux4_1 _4825_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ),
    .S0(net430),
    .S1(net421),
    .X(_2369_));
 sky130_fd_sc_hd__mux4_1 _4826_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ),
    .S0(net430),
    .S1(net421),
    .X(_2370_));
 sky130_fd_sc_hd__mux2_1 _4827_ (.A0(_2370_),
    .A1(_2369_),
    .S(net414),
    .X(_2371_));
 sky130_fd_sc_hd__mux2_1 _4828_ (.A0(_2371_),
    .A1(_2368_),
    .S(net408),
    .X(_0060_));
 sky130_fd_sc_hd__mux4_1 _4829_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ),
    .S0(net429),
    .S1(net420),
    .X(_2372_));
 sky130_fd_sc_hd__mux4_1 _4830_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ),
    .S0(net429),
    .S1(net420),
    .X(_2373_));
 sky130_fd_sc_hd__mux2_1 _4831_ (.A0(_2372_),
    .A1(_2373_),
    .S(net411),
    .X(_2374_));
 sky130_fd_sc_hd__mux4_1 _4832_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ),
    .S0(net429),
    .S1(net420),
    .X(_2375_));
 sky130_fd_sc_hd__mux4_1 _4833_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ),
    .S0(net429),
    .S1(net420),
    .X(_2376_));
 sky130_fd_sc_hd__mux2_1 _4834_ (.A0(_2376_),
    .A1(_2375_),
    .S(net414),
    .X(_2377_));
 sky130_fd_sc_hd__mux2_1 _4835_ (.A0(_2377_),
    .A1(_2374_),
    .S(net408),
    .X(_0061_));
 sky130_fd_sc_hd__mux4_1 _4836_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ),
    .S0(net429),
    .S1(net420),
    .X(_2378_));
 sky130_fd_sc_hd__mux4_1 _4837_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ),
    .S0(net429),
    .S1(net420),
    .X(_2379_));
 sky130_fd_sc_hd__mux2_1 _4838_ (.A0(_2378_),
    .A1(_2379_),
    .S(net412),
    .X(_2380_));
 sky130_fd_sc_hd__mux4_1 _4839_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ),
    .S0(net429),
    .S1(net420),
    .X(_2381_));
 sky130_fd_sc_hd__mux4_1 _4840_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ),
    .S0(net429),
    .S1(net420),
    .X(_2382_));
 sky130_fd_sc_hd__mux2_1 _4841_ (.A0(_2382_),
    .A1(_2381_),
    .S(net412),
    .X(_2383_));
 sky130_fd_sc_hd__mux2_1 _4842_ (.A0(_2383_),
    .A1(_2380_),
    .S(net407),
    .X(_0062_));
 sky130_fd_sc_hd__mux4_1 _4843_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ),
    .S0(net434),
    .S1(net423),
    .X(_2384_));
 sky130_fd_sc_hd__mux4_1 _4844_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ),
    .S0(net433),
    .S1(net423),
    .X(_2385_));
 sky130_fd_sc_hd__mux2_1 _4845_ (.A0(_2384_),
    .A1(_2385_),
    .S(net413),
    .X(_2386_));
 sky130_fd_sc_hd__mux4_1 _4846_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ),
    .S0(net433),
    .S1(net424),
    .X(_2387_));
 sky130_fd_sc_hd__mux4_1 _4847_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ),
    .S0(net433),
    .S1(net423),
    .X(_2388_));
 sky130_fd_sc_hd__mux2_1 _4848_ (.A0(_2388_),
    .A1(_2387_),
    .S(net413),
    .X(_2389_));
 sky130_fd_sc_hd__mux2_1 _4849_ (.A0(_2389_),
    .A1(_2386_),
    .S(net408),
    .X(_0063_));
 sky130_fd_sc_hd__mux4_1 _4850_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ),
    .S0(net431),
    .S1(net422),
    .X(_2390_));
 sky130_fd_sc_hd__mux4_1 _4851_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ),
    .S0(net429),
    .S1(net420),
    .X(_2391_));
 sky130_fd_sc_hd__mux2_1 _4852_ (.A0(_2390_),
    .A1(_2391_),
    .S(net412),
    .X(_2392_));
 sky130_fd_sc_hd__mux4_1 _4853_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ),
    .S0(net429),
    .S1(net420),
    .X(_2393_));
 sky130_fd_sc_hd__mux4_1 _4854_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ),
    .S0(net429),
    .S1(net420),
    .X(_2394_));
 sky130_fd_sc_hd__mux2_1 _4855_ (.A0(_2394_),
    .A1(_2393_),
    .S(net412),
    .X(_2395_));
 sky130_fd_sc_hd__mux2_1 _4856_ (.A0(_2395_),
    .A1(_2392_),
    .S(net407),
    .X(_0033_));
 sky130_fd_sc_hd__mux4_1 _4857_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ),
    .S0(net425),
    .S1(net415),
    .X(_2396_));
 sky130_fd_sc_hd__mux4_1 _4858_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ),
    .S0(net427),
    .S1(net418),
    .X(_2397_));
 sky130_fd_sc_hd__mux2_1 _4859_ (.A0(_2396_),
    .A1(_2397_),
    .S(net410),
    .X(_2398_));
 sky130_fd_sc_hd__mux4_1 _4860_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ),
    .S0(net427),
    .S1(net418),
    .X(_2399_));
 sky130_fd_sc_hd__mux4_1 _4861_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ),
    .S0(net427),
    .S1(net418),
    .X(_2400_));
 sky130_fd_sc_hd__mux2_1 _4862_ (.A0(_2400_),
    .A1(_2399_),
    .S(net411),
    .X(_2401_));
 sky130_fd_sc_hd__mux2_1 _4863_ (.A0(_2401_),
    .A1(_2398_),
    .S(net408),
    .X(_0034_));
 sky130_fd_sc_hd__mux4_1 _4864_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ),
    .S0(net432),
    .S1(net422),
    .X(_2402_));
 sky130_fd_sc_hd__mux4_1 _4865_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ),
    .S0(net432),
    .S1(net422),
    .X(_2403_));
 sky130_fd_sc_hd__mux2_1 _4866_ (.A0(_2402_),
    .A1(_2403_),
    .S(net413),
    .X(_2404_));
 sky130_fd_sc_hd__mux4_1 _4867_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ),
    .S0(net431),
    .S1(net422),
    .X(_2405_));
 sky130_fd_sc_hd__mux4_1 _4868_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ),
    .S0(net431),
    .S1(net422),
    .X(_2406_));
 sky130_fd_sc_hd__mux2_1 _4869_ (.A0(_2406_),
    .A1(_2405_),
    .S(net412),
    .X(_2407_));
 sky130_fd_sc_hd__mux2_1 _4870_ (.A0(_2407_),
    .A1(_2404_),
    .S(net407),
    .X(_0035_));
 sky130_fd_sc_hd__mux4_1 _4871_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ),
    .S0(net427),
    .S1(net418),
    .X(_2408_));
 sky130_fd_sc_hd__mux4_1 _4872_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ),
    .S0(net427),
    .S1(net418),
    .X(_2409_));
 sky130_fd_sc_hd__mux2_1 _4873_ (.A0(_2408_),
    .A1(_2409_),
    .S(net411),
    .X(_2410_));
 sky130_fd_sc_hd__mux4_1 _4874_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ),
    .S0(net427),
    .S1(net418),
    .X(_2411_));
 sky130_fd_sc_hd__mux4_1 _4875_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ),
    .S0(net427),
    .S1(net418),
    .X(_2412_));
 sky130_fd_sc_hd__mux2_1 _4876_ (.A0(_2412_),
    .A1(_2411_),
    .S(net411),
    .X(_2413_));
 sky130_fd_sc_hd__mux2_1 _4877_ (.A0(_2413_),
    .A1(_2410_),
    .S(net408),
    .X(_0036_));
 sky130_fd_sc_hd__mux4_1 _4878_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ),
    .S0(net429),
    .S1(net420),
    .X(_2414_));
 sky130_fd_sc_hd__mux4_1 _4879_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ),
    .S0(net428),
    .S1(net419),
    .X(_2415_));
 sky130_fd_sc_hd__mux2_1 _4880_ (.A0(_2414_),
    .A1(_2415_),
    .S(net411),
    .X(_2416_));
 sky130_fd_sc_hd__mux4_1 _4881_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ),
    .S0(net429),
    .S1(net420),
    .X(_2417_));
 sky130_fd_sc_hd__mux4_1 _4882_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ),
    .S0(net429),
    .S1(net420),
    .X(_2418_));
 sky130_fd_sc_hd__mux2_1 _4883_ (.A0(_2418_),
    .A1(_2417_),
    .S(net411),
    .X(_2419_));
 sky130_fd_sc_hd__mux2_1 _4884_ (.A0(_2419_),
    .A1(_2416_),
    .S(net408),
    .X(_0037_));
 sky130_fd_sc_hd__mux4_1 _4885_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ),
    .S0(net431),
    .S1(net422),
    .X(_2420_));
 sky130_fd_sc_hd__mux4_1 _4886_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ),
    .S0(net431),
    .S1(net422),
    .X(_2421_));
 sky130_fd_sc_hd__mux2_1 _4887_ (.A0(_2420_),
    .A1(_2421_),
    .S(net412),
    .X(_2422_));
 sky130_fd_sc_hd__mux4_1 _4888_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ),
    .S0(net431),
    .S1(net422),
    .X(_2423_));
 sky130_fd_sc_hd__mux4_1 _4889_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ),
    .S0(net431),
    .S1(net422),
    .X(_2424_));
 sky130_fd_sc_hd__mux2_1 _4890_ (.A0(_2424_),
    .A1(_2423_),
    .S(net413),
    .X(_2425_));
 sky130_fd_sc_hd__mux2_1 _4891_ (.A0(_2425_),
    .A1(_2422_),
    .S(net407),
    .X(_0038_));
 sky130_fd_sc_hd__mux4_1 _4892_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ),
    .S0(net427),
    .S1(net419),
    .X(_2426_));
 sky130_fd_sc_hd__mux4_1 _4893_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ),
    .S0(net428),
    .S1(net418),
    .X(_2427_));
 sky130_fd_sc_hd__mux2_1 _4894_ (.A0(_2426_),
    .A1(_2427_),
    .S(net411),
    .X(_2428_));
 sky130_fd_sc_hd__mux4_1 _4895_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ),
    .S0(net427),
    .S1(net418),
    .X(_2429_));
 sky130_fd_sc_hd__mux4_1 _4896_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ),
    .S0(net428),
    .S1(net419),
    .X(_2430_));
 sky130_fd_sc_hd__mux2_1 _4897_ (.A0(_2430_),
    .A1(_2429_),
    .S(net411),
    .X(_2431_));
 sky130_fd_sc_hd__mux2_1 _4898_ (.A0(_2431_),
    .A1(_2428_),
    .S(net408),
    .X(_0039_));
 sky130_fd_sc_hd__mux4_1 _4899_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ),
    .S0(net426),
    .S1(net417),
    .X(_2432_));
 sky130_fd_sc_hd__mux4_1 _4900_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ),
    .S0(net426),
    .S1(net417),
    .X(_2433_));
 sky130_fd_sc_hd__mux2_1 _4901_ (.A0(_2432_),
    .A1(_2433_),
    .S(net414),
    .X(_2434_));
 sky130_fd_sc_hd__mux4_1 _4902_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ),
    .S0(net426),
    .S1(net417),
    .X(_2435_));
 sky130_fd_sc_hd__mux4_1 _4903_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ),
    .S0(net426),
    .S1(net417),
    .X(_2436_));
 sky130_fd_sc_hd__mux2_1 _4904_ (.A0(_2436_),
    .A1(_2435_),
    .S(net410),
    .X(_2437_));
 sky130_fd_sc_hd__mux2_1 _4905_ (.A0(_2437_),
    .A1(_2434_),
    .S(net409),
    .X(_0040_));
 sky130_fd_sc_hd__mux4_1 _4906_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ),
    .S0(net431),
    .S1(net422),
    .X(_2438_));
 sky130_fd_sc_hd__mux4_1 _4907_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ),
    .S0(net431),
    .S1(net422),
    .X(_2439_));
 sky130_fd_sc_hd__mux2_1 _4908_ (.A0(_2438_),
    .A1(_2439_),
    .S(net412),
    .X(_2440_));
 sky130_fd_sc_hd__mux4_1 _4909_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ),
    .S0(net433),
    .S1(net423),
    .X(_2441_));
 sky130_fd_sc_hd__mux4_1 _4910_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ),
    .S0(net433),
    .S1(net423),
    .X(_2442_));
 sky130_fd_sc_hd__mux2_1 _4911_ (.A0(_2442_),
    .A1(_2441_),
    .S(net412),
    .X(_2443_));
 sky130_fd_sc_hd__mux2_1 _4912_ (.A0(_2443_),
    .A1(_2440_),
    .S(net407),
    .X(_0041_));
 sky130_fd_sc_hd__mux4_1 _4913_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ),
    .S0(net428),
    .S1(net419),
    .X(_2444_));
 sky130_fd_sc_hd__mux4_1 _4914_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ),
    .S0(net428),
    .S1(net419),
    .X(_2445_));
 sky130_fd_sc_hd__mux2_1 _4915_ (.A0(_2444_),
    .A1(_2445_),
    .S(net411),
    .X(_2446_));
 sky130_fd_sc_hd__mux4_1 _4916_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ),
    .S0(net428),
    .S1(net419),
    .X(_2447_));
 sky130_fd_sc_hd__mux4_1 _4917_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ),
    .S0(net428),
    .S1(net419),
    .X(_2448_));
 sky130_fd_sc_hd__mux2_1 _4918_ (.A0(_2448_),
    .A1(_2447_),
    .S(net411),
    .X(_2449_));
 sky130_fd_sc_hd__mux2_1 _4919_ (.A0(_2449_),
    .A1(_2446_),
    .S(net408),
    .X(_0042_));
 sky130_fd_sc_hd__mux4_1 _4920_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ),
    .S0(net425),
    .S1(net415),
    .X(_2450_));
 sky130_fd_sc_hd__mux4_1 _4921_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ),
    .S0(net425),
    .S1(net416),
    .X(_2451_));
 sky130_fd_sc_hd__mux2_1 _4922_ (.A0(_2450_),
    .A1(_2451_),
    .S(net410),
    .X(_2452_));
 sky130_fd_sc_hd__mux4_1 _4923_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ),
    .S0(net425),
    .S1(net415),
    .X(_2453_));
 sky130_fd_sc_hd__mux4_1 _4924_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ),
    .S0(net425),
    .S1(net415),
    .X(_2454_));
 sky130_fd_sc_hd__mux2_1 _4925_ (.A0(_2454_),
    .A1(_2453_),
    .S(net410),
    .X(_2455_));
 sky130_fd_sc_hd__mux2_1 _4926_ (.A0(_2455_),
    .A1(_2452_),
    .S(net409),
    .X(_0044_));
 sky130_fd_sc_hd__mux4_1 _4927_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ),
    .S0(net426),
    .S1(net416),
    .X(_2456_));
 sky130_fd_sc_hd__mux4_1 _4928_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ),
    .S0(net426),
    .S1(net415),
    .X(_2457_));
 sky130_fd_sc_hd__mux2_1 _4929_ (.A0(_2456_),
    .A1(_2457_),
    .S(net410),
    .X(_2458_));
 sky130_fd_sc_hd__mux4_1 _4930_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ),
    .S0(net425),
    .S1(net416),
    .X(_2459_));
 sky130_fd_sc_hd__mux4_1 _4931_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ),
    .S0(net426),
    .S1(net415),
    .X(_2460_));
 sky130_fd_sc_hd__mux2_1 _4932_ (.A0(_2460_),
    .A1(_2459_),
    .S(net410),
    .X(_2461_));
 sky130_fd_sc_hd__mux2_1 _4933_ (.A0(_2461_),
    .A1(_2458_),
    .S(net409),
    .X(_0045_));
 sky130_fd_sc_hd__mux4_1 _4934_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ),
    .S0(net430),
    .S1(net421),
    .X(_2462_));
 sky130_fd_sc_hd__mux4_1 _4935_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ),
    .S0(net430),
    .S1(net421),
    .X(_2463_));
 sky130_fd_sc_hd__mux2_1 _4936_ (.A0(_2462_),
    .A1(_2463_),
    .S(net411),
    .X(_2464_));
 sky130_fd_sc_hd__mux4_1 _4937_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ),
    .S0(net427),
    .S1(net418),
    .X(_2465_));
 sky130_fd_sc_hd__mux4_1 _4938_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ),
    .S0(net430),
    .S1(net421),
    .X(_2466_));
 sky130_fd_sc_hd__mux2_1 _4939_ (.A0(_2466_),
    .A1(_2465_),
    .S(net411),
    .X(_2467_));
 sky130_fd_sc_hd__mux2_1 _4940_ (.A0(_2467_),
    .A1(_2464_),
    .S(net408),
    .X(_0046_));
 sky130_fd_sc_hd__mux4_1 _4941_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ),
    .S0(net425),
    .S1(net415),
    .X(_2468_));
 sky130_fd_sc_hd__mux4_1 _4942_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ),
    .S0(net426),
    .S1(net416),
    .X(_2469_));
 sky130_fd_sc_hd__mux2_1 _4943_ (.A0(_2468_),
    .A1(_2469_),
    .S(net410),
    .X(_2470_));
 sky130_fd_sc_hd__mux4_1 _4944_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ),
    .S0(net425),
    .S1(net415),
    .X(_2471_));
 sky130_fd_sc_hd__mux4_1 _4945_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ),
    .S0(net425),
    .S1(net415),
    .X(_2472_));
 sky130_fd_sc_hd__mux2_1 _4946_ (.A0(_2472_),
    .A1(_2471_),
    .S(net410),
    .X(_2473_));
 sky130_fd_sc_hd__mux2_1 _4947_ (.A0(_2473_),
    .A1(_2470_),
    .S(net409),
    .X(_0047_));
 sky130_fd_sc_hd__mux4_1 _4948_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ),
    .S0(net433),
    .S1(net424),
    .X(_2474_));
 sky130_fd_sc_hd__mux4_1 _4949_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ),
    .S0(net433),
    .S1(net423),
    .X(_2475_));
 sky130_fd_sc_hd__mux2_1 _4950_ (.A0(_2474_),
    .A1(_2475_),
    .S(net413),
    .X(_2476_));
 sky130_fd_sc_hd__mux4_1 _4951_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ),
    .S0(net431),
    .S1(net424),
    .X(_2477_));
 sky130_fd_sc_hd__mux4_1 _4952_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ),
    .S0(net433),
    .S1(net423),
    .X(_2478_));
 sky130_fd_sc_hd__mux2_1 _4953_ (.A0(_2478_),
    .A1(_2477_),
    .S(net413),
    .X(_2479_));
 sky130_fd_sc_hd__mux2_1 _4954_ (.A0(_2479_),
    .A1(_2476_),
    .S(net407),
    .X(_0048_));
 sky130_fd_sc_hd__mux4_1 _4955_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ),
    .S0(net425),
    .S1(net415),
    .X(_2480_));
 sky130_fd_sc_hd__mux4_1 _4956_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .S1(net416),
    .X(_2481_));
 sky130_fd_sc_hd__mux2_1 _4957_ (.A0(_2480_),
    .A1(_2481_),
    .S(net410),
    .X(_2482_));
 sky130_fd_sc_hd__mux4_1 _4958_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ),
    .S0(net425),
    .S1(net415),
    .X(_2483_));
 sky130_fd_sc_hd__mux4_1 _4959_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ),
    .S0(net425),
    .S1(net415),
    .X(_2484_));
 sky130_fd_sc_hd__mux2_1 _4960_ (.A0(_2484_),
    .A1(_2483_),
    .S(net410),
    .X(_2485_));
 sky130_fd_sc_hd__mux2_1 _4961_ (.A0(_2485_),
    .A1(_2482_),
    .S(net409),
    .X(_0049_));
 sky130_fd_sc_hd__mux4_1 _4962_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ),
    .S0(net426),
    .S1(net416),
    .X(_2486_));
 sky130_fd_sc_hd__mux4_1 _4963_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .S1(net416),
    .X(_2487_));
 sky130_fd_sc_hd__mux2_1 _4964_ (.A0(_2486_),
    .A1(_2487_),
    .S(net414),
    .X(_2488_));
 sky130_fd_sc_hd__mux4_1 _4965_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ),
    .S0(net425),
    .S1(net415),
    .X(_2489_));
 sky130_fd_sc_hd__mux4_1 _4966_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ),
    .S0(net425),
    .S1(net415),
    .X(_2490_));
 sky130_fd_sc_hd__mux2_1 _4967_ (.A0(_2490_),
    .A1(_2489_),
    .S(net410),
    .X(_2491_));
 sky130_fd_sc_hd__mux2_1 _4968_ (.A0(_2491_),
    .A1(_2488_),
    .S(net409),
    .X(_0050_));
 sky130_fd_sc_hd__mux4_1 _4969_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ),
    .S0(net434),
    .S1(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ),
    .X(_2492_));
 sky130_fd_sc_hd__mux4_1 _4970_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ),
    .S0(net427),
    .S1(net418),
    .X(_2493_));
 sky130_fd_sc_hd__mux2_1 _4971_ (.A0(_2492_),
    .A1(_2493_),
    .S(net414),
    .X(_2494_));
 sky130_fd_sc_hd__mux4_1 _4972_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ),
    .S0(net434),
    .S1(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ),
    .X(_2495_));
 sky130_fd_sc_hd__mux4_1 _4973_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ),
    .S0(net427),
    .S1(net418),
    .X(_2496_));
 sky130_fd_sc_hd__mux2_1 _4974_ (.A0(_2496_),
    .A1(_2495_),
    .S(net414),
    .X(_2497_));
 sky130_fd_sc_hd__mux2_1 _4975_ (.A0(_2497_),
    .A1(_2494_),
    .S(net408),
    .X(_0051_));
 sky130_fd_sc_hd__mux4_1 _4976_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ),
    .S0(net425),
    .S1(net415),
    .X(_2498_));
 sky130_fd_sc_hd__mux4_1 _4977_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ),
    .S0(net425),
    .S1(net416),
    .X(_2499_));
 sky130_fd_sc_hd__mux2_1 _4978_ (.A0(_2498_),
    .A1(_2499_),
    .S(net410),
    .X(_2500_));
 sky130_fd_sc_hd__mux4_1 _4979_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ),
    .S0(net426),
    .S1(net417),
    .X(_2501_));
 sky130_fd_sc_hd__mux4_1 _4980_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ),
    .S0(net426),
    .S1(net417),
    .X(_2502_));
 sky130_fd_sc_hd__mux2_1 _4981_ (.A0(_2502_),
    .A1(_2501_),
    .S(net410),
    .X(_2503_));
 sky130_fd_sc_hd__mux2_1 _4982_ (.A0(_2503_),
    .A1(_2500_),
    .S(net409),
    .X(_0052_));
 sky130_fd_sc_hd__mux4_1 _4983_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ),
    .S0(net426),
    .S1(net417),
    .X(_2504_));
 sky130_fd_sc_hd__mux4_1 _4984_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ),
    .S0(net426),
    .S1(net417),
    .X(_2505_));
 sky130_fd_sc_hd__mux2_1 _4985_ (.A0(_2504_),
    .A1(_2505_),
    .S(net410),
    .X(_2506_));
 sky130_fd_sc_hd__mux4_1 _4986_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ),
    .S0(net426),
    .S1(net417),
    .X(_2507_));
 sky130_fd_sc_hd__mux4_1 _4987_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ),
    .S0(net426),
    .S1(net417),
    .X(_2508_));
 sky130_fd_sc_hd__mux2_1 _4988_ (.A0(_2508_),
    .A1(_2507_),
    .S(net410),
    .X(_2509_));
 sky130_fd_sc_hd__mux2_1 _4989_ (.A0(_2509_),
    .A1(_2506_),
    .S(net409),
    .X(_0053_));
 sky130_fd_sc_hd__mux4_1 _4990_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ),
    .S0(net432),
    .S1(net424),
    .X(_2510_));
 sky130_fd_sc_hd__mux4_1 _4991_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ),
    .S0(net432),
    .S1(net424),
    .X(_2511_));
 sky130_fd_sc_hd__mux2_1 _4992_ (.A0(_2510_),
    .A1(_2511_),
    .S(net413),
    .X(_2512_));
 sky130_fd_sc_hd__mux4_1 _4993_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ),
    .S0(net432),
    .S1(net424),
    .X(_2513_));
 sky130_fd_sc_hd__mux4_1 _4994_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ),
    .S0(net432),
    .S1(net424),
    .X(_2514_));
 sky130_fd_sc_hd__mux2_1 _4995_ (.A0(_2514_),
    .A1(_2513_),
    .S(net413),
    .X(_2515_));
 sky130_fd_sc_hd__mux2_1 _4996_ (.A0(_2515_),
    .A1(_2512_),
    .S(net407),
    .X(_0055_));
 sky130_fd_sc_hd__mux4_1 _4997_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ),
    .S0(net427),
    .S1(net418),
    .X(_2516_));
 sky130_fd_sc_hd__mux4_1 _4998_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ),
    .S0(net427),
    .S1(net418),
    .X(_2517_));
 sky130_fd_sc_hd__mux2_1 _4999_ (.A0(_2516_),
    .A1(_2517_),
    .S(net410),
    .X(_2518_));
 sky130_fd_sc_hd__mux4_1 _5000_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ),
    .S0(net427),
    .S1(net418),
    .X(_2519_));
 sky130_fd_sc_hd__mux4_1 _5001_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ),
    .S0(net427),
    .S1(net418),
    .X(_2520_));
 sky130_fd_sc_hd__mux2_1 _5002_ (.A0(_2520_),
    .A1(_2519_),
    .S(net414),
    .X(_2521_));
 sky130_fd_sc_hd__mux2_1 _5003_ (.A0(_2521_),
    .A1(_2518_),
    .S(net408),
    .X(_0056_));
 sky130_fd_sc_hd__and2_1 _5004_ (.A(net443),
    .B(net634),
    .X(_0193_));
 sky130_fd_sc_hd__and2_1 _5005_ (.A(net443),
    .B(net671),
    .X(_0194_));
 sky130_fd_sc_hd__and2_4 _5006_ (.A(net463),
    .B(net180),
    .X(_2522_));
 sky130_fd_sc_hd__mux2_1 _5007_ (.A0(net2100),
    .A1(net1117),
    .S(net295),
    .X(_2523_));
 sky130_fd_sc_hd__or3b_1 _5008_ (.A(net466),
    .B(_2523_),
    .C_N(net2085),
    .X(_0225_));
 sky130_fd_sc_hd__or2_1 _5009_ (.A(net894),
    .B(net281),
    .X(_2524_));
 sky130_fd_sc_hd__o211a_1 _5010_ (.A1(net2004),
    .A2(net298),
    .B1(net168),
    .C1(_2524_),
    .X(_0226_));
 sky130_fd_sc_hd__or2_1 _5011_ (.A(net838),
    .B(net287),
    .X(_2525_));
 sky130_fd_sc_hd__o211a_1 _5012_ (.A1(net2054),
    .A2(net300),
    .B1(net170),
    .C1(_2525_),
    .X(_0227_));
 sky130_fd_sc_hd__or2_1 _5013_ (.A(net886),
    .B(net281),
    .X(_2526_));
 sky130_fd_sc_hd__o211a_1 _5014_ (.A1(net1993),
    .A2(net298),
    .B1(net169),
    .C1(_2526_),
    .X(_0228_));
 sky130_fd_sc_hd__or2_1 _5015_ (.A(net882),
    .B(net282),
    .X(_2527_));
 sky130_fd_sc_hd__o211a_1 _5016_ (.A1(net1992),
    .A2(net298),
    .B1(net168),
    .C1(_2527_),
    .X(_0229_));
 sky130_fd_sc_hd__or2_1 _5017_ (.A(net930),
    .B(net287),
    .X(_2528_));
 sky130_fd_sc_hd__o211a_1 _5018_ (.A1(net2017),
    .A2(net300),
    .B1(net170),
    .C1(_2528_),
    .X(_0230_));
 sky130_fd_sc_hd__or2_1 _5019_ (.A(net762),
    .B(net287),
    .X(_2529_));
 sky130_fd_sc_hd__o211a_1 _5020_ (.A1(net2061),
    .A2(net300),
    .B1(net170),
    .C1(_2529_),
    .X(_0231_));
 sky130_fd_sc_hd__or2_1 _5021_ (.A(net919),
    .B(net288),
    .X(_2530_));
 sky130_fd_sc_hd__o211a_1 _5022_ (.A1(net2013),
    .A2(net300),
    .B1(net170),
    .C1(_2530_),
    .X(_0232_));
 sky130_fd_sc_hd__or2_1 _5023_ (.A(net901),
    .B(net282),
    .X(_2531_));
 sky130_fd_sc_hd__o211a_1 _5024_ (.A1(net2044),
    .A2(net298),
    .B1(net169),
    .C1(_2531_),
    .X(_0233_));
 sky130_fd_sc_hd__or2_1 _5025_ (.A(net832),
    .B(net279),
    .X(_2532_));
 sky130_fd_sc_hd__o211a_1 _5026_ (.A1(net2060),
    .A2(net297),
    .B1(net168),
    .C1(_2532_),
    .X(_0234_));
 sky130_fd_sc_hd__or2_1 _5027_ (.A(net834),
    .B(net287),
    .X(_2533_));
 sky130_fd_sc_hd__o211a_1 _5028_ (.A1(net2027),
    .A2(net300),
    .B1(net170),
    .C1(_2533_),
    .X(_0235_));
 sky130_fd_sc_hd__or2_1 _5029_ (.A(net807),
    .B(net279),
    .X(_2534_));
 sky130_fd_sc_hd__o211a_1 _5030_ (.A1(net1971),
    .A2(net297),
    .B1(net168),
    .C1(_2534_),
    .X(_0236_));
 sky130_fd_sc_hd__or2_1 _5031_ (.A(net1041),
    .B(net279),
    .X(_2535_));
 sky130_fd_sc_hd__o211a_1 _5032_ (.A1(net1989),
    .A2(net297),
    .B1(net168),
    .C1(_2535_),
    .X(_0237_));
 sky130_fd_sc_hd__or2_1 _5033_ (.A(net856),
    .B(net279),
    .X(_2536_));
 sky130_fd_sc_hd__o211a_1 _5034_ (.A1(net2015),
    .A2(net297),
    .B1(net168),
    .C1(_2536_),
    .X(_0238_));
 sky130_fd_sc_hd__or2_1 _5035_ (.A(net1029),
    .B(net285),
    .X(_2537_));
 sky130_fd_sc_hd__o211a_1 _5036_ (.A1(net2023),
    .A2(net299),
    .B1(net169),
    .C1(_2537_),
    .X(_0239_));
 sky130_fd_sc_hd__or2_1 _5037_ (.A(net608),
    .B(net280),
    .X(_2538_));
 sky130_fd_sc_hd__o211a_1 _5038_ (.A1(net2068),
    .A2(net298),
    .B1(net168),
    .C1(_2538_),
    .X(_0240_));
 sky130_fd_sc_hd__or2_1 _5039_ (.A(net1031),
    .B(net285),
    .X(_2539_));
 sky130_fd_sc_hd__o211a_1 _5040_ (.A1(net2070),
    .A2(net299),
    .B1(net169),
    .C1(_2539_),
    .X(_0241_));
 sky130_fd_sc_hd__or2_1 _5041_ (.A(net799),
    .B(net284),
    .X(_2540_));
 sky130_fd_sc_hd__o211a_1 _5042_ (.A1(net2024),
    .A2(net299),
    .B1(net169),
    .C1(_2540_),
    .X(_0242_));
 sky130_fd_sc_hd__or2_1 _5043_ (.A(net1125),
    .B(net275),
    .X(_2541_));
 sky130_fd_sc_hd__o211a_1 _5044_ (.A1(net2064),
    .A2(net294),
    .B1(net164),
    .C1(_2541_),
    .X(_0243_));
 sky130_fd_sc_hd__or2_1 _5045_ (.A(net871),
    .B(net274),
    .X(_2542_));
 sky130_fd_sc_hd__o211a_1 _5046_ (.A1(net1874),
    .A2(net294),
    .B1(net165),
    .C1(_2542_),
    .X(_0244_));
 sky130_fd_sc_hd__or2_1 _5047_ (.A(net948),
    .B(net275),
    .X(_2543_));
 sky130_fd_sc_hd__o211a_1 _5048_ (.A1(net1988),
    .A2(net294),
    .B1(net165),
    .C1(_2543_),
    .X(_0245_));
 sky130_fd_sc_hd__or2_1 _5049_ (.A(net915),
    .B(net274),
    .X(_2544_));
 sky130_fd_sc_hd__o211a_1 _5050_ (.A1(net2021),
    .A2(net294),
    .B1(net165),
    .C1(_2544_),
    .X(_0246_));
 sky130_fd_sc_hd__or2_1 _5051_ (.A(net820),
    .B(net275),
    .X(_2545_));
 sky130_fd_sc_hd__o211a_1 _5052_ (.A1(net2059),
    .A2(net294),
    .B1(net165),
    .C1(_2545_),
    .X(_0247_));
 sky130_fd_sc_hd__or2_1 _5053_ (.A(net774),
    .B(net273),
    .X(_2546_));
 sky130_fd_sc_hd__o211a_1 _5054_ (.A1(net2055),
    .A2(net292),
    .B1(net164),
    .C1(_2546_),
    .X(_0248_));
 sky130_fd_sc_hd__or2_1 _5055_ (.A(net764),
    .B(net273),
    .X(_2547_));
 sky130_fd_sc_hd__o211a_1 _5056_ (.A1(net2052),
    .A2(net293),
    .B1(net164),
    .C1(_2547_),
    .X(_0249_));
 sky130_fd_sc_hd__or2_1 _5057_ (.A(net803),
    .B(net273),
    .X(_2548_));
 sky130_fd_sc_hd__o211a_1 _5058_ (.A1(net2029),
    .A2(net293),
    .B1(net164),
    .C1(_2548_),
    .X(_0250_));
 sky130_fd_sc_hd__or2_1 _5059_ (.A(net983),
    .B(net276),
    .X(_2549_));
 sky130_fd_sc_hd__o211a_1 _5060_ (.A1(net1954),
    .A2(net295),
    .B1(net166),
    .C1(_2549_),
    .X(_0251_));
 sky130_fd_sc_hd__or2_1 _5061_ (.A(net658),
    .B(net271),
    .X(_2550_));
 sky130_fd_sc_hd__o211a_1 _5062_ (.A1(net2031),
    .A2(net292),
    .B1(net164),
    .C1(_2550_),
    .X(_0252_));
 sky130_fd_sc_hd__or2_1 _5063_ (.A(net1281),
    .B(net271),
    .X(_2551_));
 sky130_fd_sc_hd__o211a_1 _5064_ (.A1(net1887),
    .A2(net292),
    .B1(net164),
    .C1(_2551_),
    .X(_0253_));
 sky130_fd_sc_hd__or2_1 _5065_ (.A(net772),
    .B(net271),
    .X(_2552_));
 sky130_fd_sc_hd__o211a_1 _5066_ (.A1(net2036),
    .A2(net292),
    .B1(net164),
    .C1(_2552_),
    .X(_0254_));
 sky130_fd_sc_hd__nand2_1 _5067_ (.A(_1278_),
    .B(net296),
    .Y(_2553_));
 sky130_fd_sc_hd__o211a_1 _5068_ (.A1(net21),
    .A2(net296),
    .B1(net167),
    .C1(_2553_),
    .X(_0255_));
 sky130_fd_sc_hd__or2_1 _5069_ (.A(net2048),
    .B(net279),
    .X(_2554_));
 sky130_fd_sc_hd__o211a_1 _5070_ (.A1(net24),
    .A2(net297),
    .B1(net168),
    .C1(_2554_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5071_ (.A0(net25),
    .A1(net2071),
    .S(net296),
    .X(_2555_));
 sky130_fd_sc_hd__or3b_1 _5072_ (.A(net468),
    .B(_2555_),
    .C_N(net175),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5073_ (.A0(net26),
    .A1(net2144),
    .S(net296),
    .X(_2556_));
 sky130_fd_sc_hd__or3b_1 _5074_ (.A(net468),
    .B(_2556_),
    .C_N(net175),
    .X(_0258_));
 sky130_fd_sc_hd__nand2_1 _5075_ (.A(_1277_),
    .B(net296),
    .Y(_2557_));
 sky130_fd_sc_hd__o211a_1 _5076_ (.A1(net27),
    .A2(net296),
    .B1(net167),
    .C1(_2557_),
    .X(_0259_));
 sky130_fd_sc_hd__or2_1 _5077_ (.A(net877),
    .B(net289),
    .X(_2558_));
 sky130_fd_sc_hd__o211a_1 _5078_ (.A1(net28),
    .A2(net300),
    .B1(net170),
    .C1(_2558_),
    .X(_0260_));
 sky130_fd_sc_hd__or2_1 _5079_ (.A(net2151),
    .B(net279),
    .X(_2559_));
 sky130_fd_sc_hd__o211a_1 _5080_ (.A1(net29),
    .A2(net297),
    .B1(net168),
    .C1(_2559_),
    .X(_0261_));
 sky130_fd_sc_hd__or2_1 _5081_ (.A(net2153),
    .B(net290),
    .X(_2560_));
 sky130_fd_sc_hd__o211a_1 _5082_ (.A1(net30),
    .A2(net301),
    .B1(net170),
    .C1(_2560_),
    .X(_0262_));
 sky130_fd_sc_hd__or2_1 _5083_ (.A(net2107),
    .B(net289),
    .X(_2561_));
 sky130_fd_sc_hd__o211a_1 _5084_ (.A1(net1),
    .A2(net300),
    .B1(net170),
    .C1(_2561_),
    .X(_0263_));
 sky130_fd_sc_hd__or2_1 _5085_ (.A(net2131),
    .B(net277),
    .X(_2562_));
 sky130_fd_sc_hd__o211a_1 _5086_ (.A1(net2),
    .A2(net296),
    .B1(net167),
    .C1(_2562_),
    .X(_0264_));
 sky130_fd_sc_hd__or2_1 _5087_ (.A(net1698),
    .B(net276),
    .X(_2563_));
 sky130_fd_sc_hd__o211a_1 _5088_ (.A1(net3),
    .A2(net295),
    .B1(net166),
    .C1(_2563_),
    .X(_0265_));
 sky130_fd_sc_hd__or2_1 _5089_ (.A(net1998),
    .B(net289),
    .X(_2564_));
 sky130_fd_sc_hd__o211a_1 _5090_ (.A1(net4),
    .A2(net300),
    .B1(net170),
    .C1(_2564_),
    .X(_0266_));
 sky130_fd_sc_hd__or2_1 _5091_ (.A(net1990),
    .B(net289),
    .X(_2565_));
 sky130_fd_sc_hd__o211a_1 _5092_ (.A1(net5),
    .A2(net300),
    .B1(net170),
    .C1(_2565_),
    .X(_0267_));
 sky130_fd_sc_hd__or2_1 _5093_ (.A(net431),
    .B(net289),
    .X(_2566_));
 sky130_fd_sc_hd__o211a_1 _5094_ (.A1(net6),
    .A2(net300),
    .B1(net170),
    .C1(_2566_),
    .X(_0268_));
 sky130_fd_sc_hd__or2_1 _5095_ (.A(net415),
    .B(net278),
    .X(_2567_));
 sky130_fd_sc_hd__o211a_1 _5096_ (.A1(net7),
    .A2(net296),
    .B1(net167),
    .C1(_2567_),
    .X(_0269_));
 sky130_fd_sc_hd__or2_1 _5097_ (.A(net414),
    .B(net276),
    .X(_2568_));
 sky130_fd_sc_hd__o211a_1 _5098_ (.A1(net8),
    .A2(net292),
    .B1(net164),
    .C1(_2568_),
    .X(_0270_));
 sky130_fd_sc_hd__or2_1 _5099_ (.A(net409),
    .B(net276),
    .X(_2569_));
 sky130_fd_sc_hd__o211a_1 _5100_ (.A1(net9),
    .A2(net295),
    .B1(net166),
    .C1(_2569_),
    .X(_0271_));
 sky130_fd_sc_hd__or2_1 _5101_ (.A(net2126),
    .B(net284),
    .X(_2570_));
 sky130_fd_sc_hd__o211a_1 _5102_ (.A1(net10),
    .A2(net299),
    .B1(net169),
    .C1(_2570_),
    .X(_0272_));
 sky130_fd_sc_hd__or2_1 _5103_ (.A(net405),
    .B(net290),
    .X(_2571_));
 sky130_fd_sc_hd__o211a_1 _5104_ (.A1(net11),
    .A2(net301),
    .B1(_2522_),
    .C1(_2571_),
    .X(_0273_));
 sky130_fd_sc_hd__or2_1 _5105_ (.A(net386),
    .B(net278),
    .X(_2572_));
 sky130_fd_sc_hd__o211a_1 _5106_ (.A1(net12),
    .A2(net296),
    .B1(net167),
    .C1(_2572_),
    .X(_0274_));
 sky130_fd_sc_hd__or2_1 _5107_ (.A(net384),
    .B(net290),
    .X(_2573_));
 sky130_fd_sc_hd__o211a_1 _5108_ (.A1(net13),
    .A2(net301),
    .B1(_2522_),
    .C1(_2573_),
    .X(_0275_));
 sky130_fd_sc_hd__or2_1 _5109_ (.A(net380),
    .B(net275),
    .X(_2574_));
 sky130_fd_sc_hd__o211a_1 _5110_ (.A1(net14),
    .A2(net294),
    .B1(net165),
    .C1(_2574_),
    .X(_0276_));
 sky130_fd_sc_hd__or2_1 _5111_ (.A(net2110),
    .B(net286),
    .X(_2575_));
 sky130_fd_sc_hd__o211a_1 _5112_ (.A1(net15),
    .A2(net299),
    .B1(net169),
    .C1(_2575_),
    .X(_0277_));
 sky130_fd_sc_hd__or2_1 _5113_ (.A(net2018),
    .B(net277),
    .X(_2576_));
 sky130_fd_sc_hd__o211a_1 _5114_ (.A1(net16),
    .A2(net296),
    .B1(net167),
    .C1(_2576_),
    .X(_0278_));
 sky130_fd_sc_hd__or2_1 _5115_ (.A(net1972),
    .B(net276),
    .X(_2577_));
 sky130_fd_sc_hd__o211a_1 _5116_ (.A1(net17),
    .A2(net295),
    .B1(net166),
    .C1(_2577_),
    .X(_0279_));
 sky130_fd_sc_hd__or2_1 _5117_ (.A(net2116),
    .B(net286),
    .X(_2578_));
 sky130_fd_sc_hd__o211a_1 _5118_ (.A1(net18),
    .A2(net299),
    .B1(net169),
    .C1(_2578_),
    .X(_0280_));
 sky130_fd_sc_hd__or2_1 _5119_ (.A(net1742),
    .B(net276),
    .X(_2579_));
 sky130_fd_sc_hd__o211a_1 _5120_ (.A1(net19),
    .A2(net295),
    .B1(net166),
    .C1(_2579_),
    .X(_0281_));
 sky130_fd_sc_hd__or2_1 _5121_ (.A(net2073),
    .B(net289),
    .X(_2580_));
 sky130_fd_sc_hd__o211a_1 _5122_ (.A1(net20),
    .A2(net300),
    .B1(net170),
    .C1(_2580_),
    .X(_0282_));
 sky130_fd_sc_hd__or2_1 _5123_ (.A(net2091),
    .B(net273),
    .X(_2581_));
 sky130_fd_sc_hd__o211a_1 _5124_ (.A1(net22),
    .A2(net293),
    .B1(net164),
    .C1(_2581_),
    .X(_0283_));
 sky130_fd_sc_hd__or2_1 _5125_ (.A(net1945),
    .B(net277),
    .X(_2582_));
 sky130_fd_sc_hd__o211a_1 _5126_ (.A1(net23),
    .A2(net296),
    .B1(net167),
    .C1(_2582_),
    .X(_0284_));
 sky130_fd_sc_hd__or2_1 _5127_ (.A(net554),
    .B(net276),
    .X(_2583_));
 sky130_fd_sc_hd__o211a_1 _5128_ (.A1(net921),
    .A2(net295),
    .B1(net166),
    .C1(_2583_),
    .X(_0285_));
 sky130_fd_sc_hd__or2_1 _5129_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[3] ),
    .B(net281),
    .X(_2584_));
 sky130_fd_sc_hd__o211a_1 _5130_ (.A1(net711),
    .A2(net298),
    .B1(net169),
    .C1(_2584_),
    .X(_0286_));
 sky130_fd_sc_hd__or2_1 _5131_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[4] ),
    .B(net281),
    .X(_2585_));
 sky130_fd_sc_hd__o211a_1 _5132_ (.A1(net880),
    .A2(net298),
    .B1(net168),
    .C1(_2585_),
    .X(_0287_));
 sky130_fd_sc_hd__or2_1 _5133_ (.A(net725),
    .B(net282),
    .X(_2586_));
 sky130_fd_sc_hd__o211a_1 _5134_ (.A1(net865),
    .A2(net298),
    .B1(net169),
    .C1(_2586_),
    .X(_0288_));
 sky130_fd_sc_hd__or2_1 _5135_ (.A(net842),
    .B(net282),
    .X(_2587_));
 sky130_fd_sc_hd__o211a_1 _5136_ (.A1(net850),
    .A2(net297),
    .B1(net168),
    .C1(_2587_),
    .X(_0289_));
 sky130_fd_sc_hd__or2_1 _5137_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[7] ),
    .B(net282),
    .X(_2588_));
 sky130_fd_sc_hd__o211a_1 _5138_ (.A1(net824),
    .A2(net298),
    .B1(net169),
    .C1(_2588_),
    .X(_0290_));
 sky130_fd_sc_hd__or2_1 _5139_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[8] ),
    .B(net281),
    .X(_2589_));
 sky130_fd_sc_hd__o211a_1 _5140_ (.A1(net544),
    .A2(net298),
    .B1(net168),
    .C1(_2589_),
    .X(_0291_));
 sky130_fd_sc_hd__or2_1 _5141_ (.A(net788),
    .B(net287),
    .X(_2590_));
 sky130_fd_sc_hd__o211a_1 _5142_ (.A1(net958),
    .A2(net300),
    .B1(net170),
    .C1(_2590_),
    .X(_0292_));
 sky130_fd_sc_hd__or2_1 _5143_ (.A(net552),
    .B(net279),
    .X(_2591_));
 sky130_fd_sc_hd__o211a_1 _5144_ (.A1(net975),
    .A2(net297),
    .B1(net168),
    .C1(_2591_),
    .X(_0293_));
 sky130_fd_sc_hd__or2_1 _5145_ (.A(net822),
    .B(net280),
    .X(_2592_));
 sky130_fd_sc_hd__o211a_1 _5146_ (.A1(net844),
    .A2(net298),
    .B1(net168),
    .C1(_2592_),
    .X(_0294_));
 sky130_fd_sc_hd__or2_1 _5147_ (.A(net580),
    .B(net289),
    .X(_2593_));
 sky130_fd_sc_hd__o211a_1 _5148_ (.A1(net826),
    .A2(net300),
    .B1(net170),
    .C1(_2593_),
    .X(_0295_));
 sky130_fd_sc_hd__or2_1 _5149_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[13] ),
    .B(net284),
    .X(_2594_));
 sky130_fd_sc_hd__o211a_1 _5150_ (.A1(net782),
    .A2(net299),
    .B1(net169),
    .C1(_2594_),
    .X(_0296_));
 sky130_fd_sc_hd__or2_1 _5151_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[14] ),
    .B(net279),
    .X(_2595_));
 sky130_fd_sc_hd__o211a_1 _5152_ (.A1(net830),
    .A2(net297),
    .B1(net168),
    .C1(_2595_),
    .X(_0297_));
 sky130_fd_sc_hd__or2_1 _5153_ (.A(net792),
    .B(net287),
    .X(_2596_));
 sky130_fd_sc_hd__o211a_1 _5154_ (.A1(net890),
    .A2(net300),
    .B1(net170),
    .C1(_2596_),
    .X(_0298_));
 sky130_fd_sc_hd__or2_1 _5155_ (.A(net548),
    .B(net283),
    .X(_2597_));
 sky130_fd_sc_hd__o211a_1 _5156_ (.A1(net816),
    .A2(net298),
    .B1(net168),
    .C1(_2597_),
    .X(_0299_));
 sky130_fd_sc_hd__or2_1 _5157_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[17] ),
    .B(net285),
    .X(_2598_));
 sky130_fd_sc_hd__o211a_1 _5158_ (.A1(net971),
    .A2(net299),
    .B1(net169),
    .C1(_2598_),
    .X(_0300_));
 sky130_fd_sc_hd__or2_1 _5159_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[18] ),
    .B(net287),
    .X(_2599_));
 sky130_fd_sc_hd__o211a_1 _5160_ (.A1(net858),
    .A2(net300),
    .B1(net170),
    .C1(_2599_),
    .X(_0301_));
 sky130_fd_sc_hd__or2_1 _5161_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[19] ),
    .B(net284),
    .X(_2600_));
 sky130_fd_sc_hd__o211a_1 _5162_ (.A1(net646),
    .A2(net299),
    .B1(net169),
    .C1(_2600_),
    .X(_0302_));
 sky130_fd_sc_hd__or2_1 _5163_ (.A(net848),
    .B(net271),
    .X(_2601_));
 sky130_fd_sc_hd__o211a_1 _5164_ (.A1(net888),
    .A2(net292),
    .B1(net164),
    .C1(_2601_),
    .X(_0303_));
 sky130_fd_sc_hd__or2_1 _5165_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[21] ),
    .B(net274),
    .X(_2602_));
 sky130_fd_sc_hd__o211a_1 _5166_ (.A1(net861),
    .A2(net294),
    .B1(net165),
    .C1(_2602_),
    .X(_0304_));
 sky130_fd_sc_hd__or2_1 _5167_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[22] ),
    .B(net275),
    .X(_2603_));
 sky130_fd_sc_hd__o211a_1 _5168_ (.A1(net854),
    .A2(net294),
    .B1(net165),
    .C1(_2603_),
    .X(_0305_));
 sky130_fd_sc_hd__or2_1 _5169_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[23] ),
    .B(net271),
    .X(_2604_));
 sky130_fd_sc_hd__o211a_1 _5170_ (.A1(net776),
    .A2(net292),
    .B1(net164),
    .C1(_2604_),
    .X(_0306_));
 sky130_fd_sc_hd__or2_1 _5171_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[24] ),
    .B(net274),
    .X(_2605_));
 sky130_fd_sc_hd__o211a_1 _5172_ (.A1(net760),
    .A2(net294),
    .B1(net165),
    .C1(_2605_),
    .X(_0307_));
 sky130_fd_sc_hd__or2_1 _5173_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[25] ),
    .B(net272),
    .X(_2606_));
 sky130_fd_sc_hd__o211a_1 _5174_ (.A1(net946),
    .A2(net292),
    .B1(net164),
    .C1(_2606_),
    .X(_0308_));
 sky130_fd_sc_hd__or2_1 _5175_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[26] ),
    .B(net274),
    .X(_2607_));
 sky130_fd_sc_hd__o211a_1 _5176_ (.A1(net896),
    .A2(net294),
    .B1(net165),
    .C1(_2607_),
    .X(_0309_));
 sky130_fd_sc_hd__or2_1 _5177_ (.A(net648),
    .B(net272),
    .X(_2608_));
 sky130_fd_sc_hd__o211a_1 _5178_ (.A1(net828),
    .A2(net293),
    .B1(net164),
    .C1(_2608_),
    .X(_0310_));
 sky130_fd_sc_hd__or2_1 _5179_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[28] ),
    .B(net271),
    .X(_2609_));
 sky130_fd_sc_hd__o211a_1 _5180_ (.A1(net846),
    .A2(net292),
    .B1(net164),
    .C1(_2609_),
    .X(_0311_));
 sky130_fd_sc_hd__or2_1 _5181_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[29] ),
    .B(net276),
    .X(_2610_));
 sky130_fd_sc_hd__o211a_1 _5182_ (.A1(net1011),
    .A2(net295),
    .B1(net166),
    .C1(_2610_),
    .X(_0312_));
 sky130_fd_sc_hd__or2_1 _5183_ (.A(net814),
    .B(net272),
    .X(_2611_));
 sky130_fd_sc_hd__o211a_1 _5184_ (.A1(net836),
    .A2(net293),
    .B1(net164),
    .C1(_2611_),
    .X(_0313_));
 sky130_fd_sc_hd__or2_1 _5185_ (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[31] ),
    .B(net272),
    .X(_2612_));
 sky130_fd_sc_hd__o211a_1 _5186_ (.A1(net818),
    .A2(net293),
    .B1(net164),
    .C1(_2612_),
    .X(_0314_));
 sky130_fd_sc_hd__or2_4 _5187_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .X(_2613_));
 sky130_fd_sc_hd__o311ai_4 _5188_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .A2(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .A3(_2613_),
    .B1(net456),
    .C1(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .Y(_2614_));
 sky130_fd_sc_hd__nand2_1 _5189_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .Y(_2615_));
 sky130_fd_sc_hd__nor2_1 _5190_ (.A(_2614_),
    .B(_2615_),
    .Y(_2616_));
 sky130_fd_sc_hd__or2_2 _5191_ (.A(_2614_),
    .B(_2615_),
    .X(_2617_));
 sky130_fd_sc_hd__and3_1 _5192_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(_1282_),
    .C(_2616_),
    .X(_2618_));
 sky130_fd_sc_hd__or3_2 _5193_ (.A(_1281_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .C(_2617_),
    .X(_2619_));
 sky130_fd_sc_hd__nor2_2 _5194_ (.A(net471),
    .B(net270),
    .Y(_2620_));
 sky130_fd_sc_hd__nand2_1 _5195_ (.A(net460),
    .B(_2619_),
    .Y(_2621_));
 sky130_fd_sc_hd__o22a_1 _5196_ (.A1(net329),
    .A2(_2619_),
    .B1(_2621_),
    .B2(net936),
    .X(_0315_));
 sky130_fd_sc_hd__a22o_1 _5197_ (.A1(net330),
    .A2(net270),
    .B1(net236),
    .B2(net1025),
    .X(_0316_));
 sky130_fd_sc_hd__o22a_1 _5198_ (.A1(net331),
    .A2(_2619_),
    .B1(_2621_),
    .B2(net995),
    .X(_0317_));
 sky130_fd_sc_hd__o22a_1 _5199_ (.A1(net332),
    .A2(_2619_),
    .B1(_2621_),
    .B2(net1724),
    .X(_0318_));
 sky130_fd_sc_hd__a22o_1 _5200_ (.A1(net327),
    .A2(net270),
    .B1(net236),
    .B2(net1073),
    .X(_0319_));
 sky130_fd_sc_hd__a22o_1 _5201_ (.A1(_1608_),
    .A2(net270),
    .B1(net236),
    .B2(net1488),
    .X(_0320_));
 sky130_fd_sc_hd__a22o_1 _5202_ (.A1(net326),
    .A2(net270),
    .B1(net236),
    .B2(net1115),
    .X(_0321_));
 sky130_fd_sc_hd__a22o_1 _5203_ (.A1(net328),
    .A2(net270),
    .B1(net236),
    .B2(net1462),
    .X(_0322_));
 sky130_fd_sc_hd__a22o_1 _5204_ (.A1(net323),
    .A2(net270),
    .B1(net236),
    .B2(net1113),
    .X(_0323_));
 sky130_fd_sc_hd__a22o_1 _5205_ (.A1(net325),
    .A2(net270),
    .B1(net236),
    .B2(net1458),
    .X(_0324_));
 sky130_fd_sc_hd__a22o_1 _5206_ (.A1(net324),
    .A2(net270),
    .B1(net236),
    .B2(net1165),
    .X(_0325_));
 sky130_fd_sc_hd__a22o_1 _5207_ (.A1(net322),
    .A2(net269),
    .B1(net235),
    .B2(net1430),
    .X(_0326_));
 sky130_fd_sc_hd__a22o_1 _5208_ (.A1(net319),
    .A2(net270),
    .B1(net236),
    .B2(net1572),
    .X(_0327_));
 sky130_fd_sc_hd__a22o_1 _5209_ (.A1(net321),
    .A2(net269),
    .B1(net235),
    .B2(net1672),
    .X(_0328_));
 sky130_fd_sc_hd__a22o_1 _5210_ (.A1(net320),
    .A2(net269),
    .B1(net235),
    .B2(net1714),
    .X(_0329_));
 sky130_fd_sc_hd__a22o_1 _5211_ (.A1(net318),
    .A2(net270),
    .B1(net236),
    .B2(net1215),
    .X(_0330_));
 sky130_fd_sc_hd__a22o_1 _5212_ (.A1(net342),
    .A2(net269),
    .B1(net235),
    .B2(net1480),
    .X(_0331_));
 sky130_fd_sc_hd__a22o_1 _5213_ (.A1(_1382_),
    .A2(net269),
    .B1(net235),
    .B2(net1099),
    .X(_0332_));
 sky130_fd_sc_hd__a22o_1 _5214_ (.A1(net341),
    .A2(net270),
    .B1(net236),
    .B2(net1351),
    .X(_0333_));
 sky130_fd_sc_hd__a22o_1 _5215_ (.A1(net343),
    .A2(net269),
    .B1(net235),
    .B2(net1119),
    .X(_0334_));
 sky130_fd_sc_hd__a22o_1 _5216_ (.A1(net338),
    .A2(net269),
    .B1(net235),
    .B2(net1516),
    .X(_0335_));
 sky130_fd_sc_hd__a22o_1 _5217_ (.A1(net340),
    .A2(net269),
    .B1(net235),
    .B2(net1133),
    .X(_0336_));
 sky130_fd_sc_hd__a22o_1 _5218_ (.A1(net339),
    .A2(net269),
    .B1(net235),
    .B2(net1596),
    .X(_0337_));
 sky130_fd_sc_hd__a22o_1 _5219_ (.A1(net337),
    .A2(net269),
    .B1(net235),
    .B2(net1167),
    .X(_0338_));
 sky130_fd_sc_hd__a22o_1 _5220_ (.A1(net334),
    .A2(net270),
    .B1(net236),
    .B2(net1496),
    .X(_0339_));
 sky130_fd_sc_hd__a22o_1 _5221_ (.A1(net336),
    .A2(net269),
    .B1(net235),
    .B2(net1546),
    .X(_0340_));
 sky130_fd_sc_hd__a22o_1 _5222_ (.A1(net335),
    .A2(net269),
    .B1(net235),
    .B2(net1129),
    .X(_0341_));
 sky130_fd_sc_hd__a22o_1 _5223_ (.A1(net333),
    .A2(net269),
    .B1(net235),
    .B2(net1464),
    .X(_0342_));
 sky130_fd_sc_hd__a22o_1 _5224_ (.A1(net346),
    .A2(net269),
    .B1(net235),
    .B2(net1093),
    .X(_0343_));
 sky130_fd_sc_hd__a22o_1 _5225_ (.A1(net344),
    .A2(net269),
    .B1(net235),
    .B2(net1612),
    .X(_0344_));
 sky130_fd_sc_hd__a22o_1 _5226_ (.A1(net345),
    .A2(net270),
    .B1(net236),
    .B2(net1736),
    .X(_0345_));
 sky130_fd_sc_hd__a22o_1 _5227_ (.A1(net368),
    .A2(net269),
    .B1(net235),
    .B2(net965),
    .X(_0346_));
 sky130_fd_sc_hd__or3_2 _5228_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(_1282_),
    .C(_2614_),
    .X(_2622_));
 sky130_fd_sc_hd__nand2_1 _5229_ (.A(_1283_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .Y(_2623_));
 sky130_fd_sc_hd__nor2_1 _5230_ (.A(_2622_),
    .B(_2623_),
    .Y(_2624_));
 sky130_fd_sc_hd__or2_1 _5231_ (.A(_2622_),
    .B(_2623_),
    .X(_2625_));
 sky130_fd_sc_hd__nor2_2 _5232_ (.A(net471),
    .B(net267),
    .Y(_2626_));
 sky130_fd_sc_hd__nand2_1 _5233_ (.A(net462),
    .B(_2625_),
    .Y(_2627_));
 sky130_fd_sc_hd__a22o_1 _5234_ (.A1(net329),
    .A2(net267),
    .B1(net234),
    .B2(net1520),
    .X(_0347_));
 sky130_fd_sc_hd__o22a_1 _5235_ (.A1(net330),
    .A2(_2625_),
    .B1(_2627_),
    .B2(net1047),
    .X(_0348_));
 sky130_fd_sc_hd__a22o_1 _5236_ (.A1(net331),
    .A2(net267),
    .B1(net234),
    .B2(net1381),
    .X(_0349_));
 sky130_fd_sc_hd__o22a_1 _5237_ (.A1(net332),
    .A2(_2625_),
    .B1(_2627_),
    .B2(net869),
    .X(_0350_));
 sky130_fd_sc_hd__a22o_1 _5238_ (.A1(net327),
    .A2(net267),
    .B1(net233),
    .B2(net1101),
    .X(_0351_));
 sky130_fd_sc_hd__a22o_1 _5239_ (.A1(_1608_),
    .A2(net267),
    .B1(net233),
    .B2(net1015),
    .X(_0352_));
 sky130_fd_sc_hd__a22o_1 _5240_ (.A1(net326),
    .A2(net267),
    .B1(net234),
    .B2(net1235),
    .X(_0353_));
 sky130_fd_sc_hd__a22o_1 _5241_ (.A1(net328),
    .A2(net267),
    .B1(net234),
    .B2(net1446),
    .X(_0354_));
 sky130_fd_sc_hd__a22o_1 _5242_ (.A1(net323),
    .A2(net267),
    .B1(net234),
    .B2(net1057),
    .X(_0355_));
 sky130_fd_sc_hd__a22o_1 _5243_ (.A1(net325),
    .A2(net267),
    .B1(net234),
    .B2(net1239),
    .X(_0356_));
 sky130_fd_sc_hd__a22o_1 _5244_ (.A1(net324),
    .A2(net268),
    .B1(net234),
    .B2(net1169),
    .X(_0357_));
 sky130_fd_sc_hd__a22o_1 _5245_ (.A1(net322),
    .A2(net268),
    .B1(net233),
    .B2(net1692),
    .X(_0358_));
 sky130_fd_sc_hd__a22o_1 _5246_ (.A1(net319),
    .A2(net267),
    .B1(net234),
    .B2(net1231),
    .X(_0359_));
 sky130_fd_sc_hd__a22o_1 _5247_ (.A1(net321),
    .A2(net268),
    .B1(net233),
    .B2(net1558),
    .X(_0360_));
 sky130_fd_sc_hd__a22o_1 _5248_ (.A1(_1679_),
    .A2(net267),
    .B1(net234),
    .B2(net1317),
    .X(_0361_));
 sky130_fd_sc_hd__a22o_1 _5249_ (.A1(net318),
    .A2(net267),
    .B1(net234),
    .B2(net1638),
    .X(_0362_));
 sky130_fd_sc_hd__a22o_1 _5250_ (.A1(net342),
    .A2(net268),
    .B1(net233),
    .B2(net1357),
    .X(_0363_));
 sky130_fd_sc_hd__a22o_1 _5251_ (.A1(_1382_),
    .A2(net268),
    .B1(net233),
    .B2(net967),
    .X(_0364_));
 sky130_fd_sc_hd__a22o_1 _5252_ (.A1(net341),
    .A2(net267),
    .B1(net234),
    .B2(net1506),
    .X(_0365_));
 sky130_fd_sc_hd__a22o_1 _5253_ (.A1(net343),
    .A2(net268),
    .B1(net233),
    .B2(net925),
    .X(_0366_));
 sky130_fd_sc_hd__a22o_1 _5254_ (.A1(net338),
    .A2(net268),
    .B1(net233),
    .B2(net1361),
    .X(_0367_));
 sky130_fd_sc_hd__a22o_1 _5255_ (.A1(net340),
    .A2(net268),
    .B1(net233),
    .B2(net1347),
    .X(_0368_));
 sky130_fd_sc_hd__a22o_1 _5256_ (.A1(net339),
    .A2(net267),
    .B1(net234),
    .B2(net1055),
    .X(_0369_));
 sky130_fd_sc_hd__a22o_1 _5257_ (.A1(net337),
    .A2(net268),
    .B1(net233),
    .B2(net1151),
    .X(_0370_));
 sky130_fd_sc_hd__a22o_1 _5258_ (.A1(net334),
    .A2(net267),
    .B1(net234),
    .B2(net1039),
    .X(_0371_));
 sky130_fd_sc_hd__a22o_1 _5259_ (.A1(net336),
    .A2(net268),
    .B1(net233),
    .B2(net1107),
    .X(_0372_));
 sky130_fd_sc_hd__a22o_1 _5260_ (.A1(net335),
    .A2(net268),
    .B1(net233),
    .B2(net1353),
    .X(_0373_));
 sky130_fd_sc_hd__a22o_1 _5261_ (.A1(net333),
    .A2(net268),
    .B1(net233),
    .B2(net1580),
    .X(_0374_));
 sky130_fd_sc_hd__a22o_1 _5262_ (.A1(net346),
    .A2(net268),
    .B1(net233),
    .B2(net1023),
    .X(_0375_));
 sky130_fd_sc_hd__a22o_1 _5263_ (.A1(net344),
    .A2(net268),
    .B1(net233),
    .B2(net1193),
    .X(_0376_));
 sky130_fd_sc_hd__a22o_1 _5264_ (.A1(net345),
    .A2(net267),
    .B1(net234),
    .B2(net989),
    .X(_0377_));
 sky130_fd_sc_hd__a22o_1 _5265_ (.A1(net368),
    .A2(net268),
    .B1(net233),
    .B2(net1179),
    .X(_0378_));
 sky130_fd_sc_hd__or3_4 _5266_ (.A(_1281_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .C(_2614_),
    .X(_2628_));
 sky130_fd_sc_hd__nor2_2 _5267_ (.A(_2623_),
    .B(_2628_),
    .Y(_2629_));
 sky130_fd_sc_hd__or2_1 _5268_ (.A(_2623_),
    .B(_2628_),
    .X(_2630_));
 sky130_fd_sc_hd__nor2_2 _5269_ (.A(net471),
    .B(net265),
    .Y(_2631_));
 sky130_fd_sc_hd__nand2_1 _5270_ (.A(net460),
    .B(_2630_),
    .Y(_2632_));
 sky130_fd_sc_hd__o22a_1 _5271_ (.A1(net329),
    .A2(_2630_),
    .B1(_2632_),
    .B2(net903),
    .X(_0379_));
 sky130_fd_sc_hd__a22o_1 _5272_ (.A1(net330),
    .A2(net266),
    .B1(net232),
    .B2(net1217),
    .X(_0380_));
 sky130_fd_sc_hd__a22o_1 _5273_ (.A1(net331),
    .A2(net266),
    .B1(net232),
    .B2(net1201),
    .X(_0381_));
 sky130_fd_sc_hd__o22a_1 _5274_ (.A1(net332),
    .A2(_2630_),
    .B1(_2632_),
    .B2(net812),
    .X(_0382_));
 sky130_fd_sc_hd__a22o_1 _5275_ (.A1(net327),
    .A2(net266),
    .B1(net231),
    .B2(net1654),
    .X(_0383_));
 sky130_fd_sc_hd__a22o_1 _5276_ (.A1(_1608_),
    .A2(net266),
    .B1(net232),
    .B2(net1033),
    .X(_0384_));
 sky130_fd_sc_hd__a22o_1 _5277_ (.A1(net326),
    .A2(net266),
    .B1(net232),
    .B2(net1219),
    .X(_0385_));
 sky130_fd_sc_hd__a22o_1 _5278_ (.A1(net328),
    .A2(net266),
    .B1(net232),
    .B2(net1554),
    .X(_0386_));
 sky130_fd_sc_hd__a22o_1 _5279_ (.A1(net323),
    .A2(net266),
    .B1(net232),
    .B2(net1263),
    .X(_0387_));
 sky130_fd_sc_hd__a22o_1 _5280_ (.A1(net325),
    .A2(net266),
    .B1(net232),
    .B2(net1365),
    .X(_0388_));
 sky130_fd_sc_hd__a22o_1 _5281_ (.A1(net324),
    .A2(net266),
    .B1(net232),
    .B2(net1021),
    .X(_0389_));
 sky130_fd_sc_hd__a22o_1 _5282_ (.A1(net322),
    .A2(net265),
    .B1(net231),
    .B2(net1620),
    .X(_0390_));
 sky130_fd_sc_hd__a22o_1 _5283_ (.A1(net319),
    .A2(net266),
    .B1(net232),
    .B2(net934),
    .X(_0391_));
 sky130_fd_sc_hd__a22o_1 _5284_ (.A1(net321),
    .A2(net265),
    .B1(net231),
    .B2(net1500),
    .X(_0392_));
 sky130_fd_sc_hd__a22o_1 _5285_ (.A1(net320),
    .A2(net265),
    .B1(net231),
    .B2(net1424),
    .X(_0393_));
 sky130_fd_sc_hd__a22o_1 _5286_ (.A1(net318),
    .A2(net266),
    .B1(net232),
    .B2(net1582),
    .X(_0394_));
 sky130_fd_sc_hd__a22o_1 _5287_ (.A1(net342),
    .A2(net265),
    .B1(net231),
    .B2(net1287),
    .X(_0395_));
 sky130_fd_sc_hd__a22o_1 _5288_ (.A1(_1382_),
    .A2(net265),
    .B1(net231),
    .B2(net997),
    .X(_0396_));
 sky130_fd_sc_hd__a22o_1 _5289_ (.A1(net341),
    .A2(net266),
    .B1(net232),
    .B2(net1267),
    .X(_0397_));
 sky130_fd_sc_hd__a22o_1 _5290_ (.A1(net343),
    .A2(net265),
    .B1(net231),
    .B2(net1440),
    .X(_0398_));
 sky130_fd_sc_hd__a22o_1 _5291_ (.A1(net338),
    .A2(net265),
    .B1(net231),
    .B2(net1650),
    .X(_0399_));
 sky130_fd_sc_hd__a22o_1 _5292_ (.A1(net340),
    .A2(net265),
    .B1(net231),
    .B2(net1037),
    .X(_0400_));
 sky130_fd_sc_hd__a22o_1 _5293_ (.A1(net339),
    .A2(net266),
    .B1(net232),
    .B2(net1510),
    .X(_0401_));
 sky130_fd_sc_hd__a22o_1 _5294_ (.A1(net337),
    .A2(net265),
    .B1(net231),
    .B2(net1680),
    .X(_0402_));
 sky130_fd_sc_hd__a22o_1 _5295_ (.A1(net334),
    .A2(net266),
    .B1(net232),
    .B2(net1059),
    .X(_0403_));
 sky130_fd_sc_hd__a22o_1 _5296_ (.A1(net336),
    .A2(net265),
    .B1(net231),
    .B2(net1686),
    .X(_0404_));
 sky130_fd_sc_hd__a22o_1 _5297_ (.A1(net335),
    .A2(net265),
    .B1(net231),
    .B2(net1614),
    .X(_0405_));
 sky130_fd_sc_hd__a22o_1 _5298_ (.A1(net333),
    .A2(net265),
    .B1(net231),
    .B2(net1303),
    .X(_0406_));
 sky130_fd_sc_hd__a22o_1 _5299_ (.A1(net346),
    .A2(net265),
    .B1(net231),
    .B2(net1369),
    .X(_0407_));
 sky130_fd_sc_hd__a22o_1 _5300_ (.A1(net344),
    .A2(net265),
    .B1(net231),
    .B2(net1826),
    .X(_0408_));
 sky130_fd_sc_hd__a22o_1 _5301_ (.A1(net345),
    .A2(net266),
    .B1(net232),
    .B2(net938),
    .X(_0409_));
 sky130_fd_sc_hd__a22o_1 _5302_ (.A1(net368),
    .A2(net265),
    .B1(net231),
    .B2(net1285),
    .X(_0410_));
 sky130_fd_sc_hd__and3_1 _5303_ (.A(_1281_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .C(_2616_),
    .X(_2633_));
 sky130_fd_sc_hd__or3_2 _5304_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(_1282_),
    .C(_2617_),
    .X(_2634_));
 sky130_fd_sc_hd__nor2_2 _5305_ (.A(net471),
    .B(net264),
    .Y(_2635_));
 sky130_fd_sc_hd__nand2_1 _5306_ (.A(net460),
    .B(_2634_),
    .Y(_2636_));
 sky130_fd_sc_hd__a22o_1 _5307_ (.A1(net329),
    .A2(net264),
    .B1(net230),
    .B2(net1604),
    .X(_0411_));
 sky130_fd_sc_hd__o22a_1 _5308_ (.A1(net330),
    .A2(_2634_),
    .B1(_2636_),
    .B2(net1660),
    .X(_0412_));
 sky130_fd_sc_hd__o22a_1 _5309_ (.A1(net331),
    .A2(_2634_),
    .B1(_2636_),
    .B2(net801),
    .X(_0413_));
 sky130_fd_sc_hd__o22a_1 _5310_ (.A1(net332),
    .A2(_2634_),
    .B1(_2636_),
    .B2(net913),
    .X(_0414_));
 sky130_fd_sc_hd__a22o_1 _5311_ (.A1(net327),
    .A2(net264),
    .B1(net230),
    .B2(net1003),
    .X(_0415_));
 sky130_fd_sc_hd__a22o_1 _5312_ (.A1(_1608_),
    .A2(net264),
    .B1(net230),
    .B2(net1502),
    .X(_0416_));
 sky130_fd_sc_hd__a22o_1 _5313_ (.A1(net326),
    .A2(net264),
    .B1(net230),
    .B2(net1478),
    .X(_0417_));
 sky130_fd_sc_hd__a22o_1 _5314_ (.A1(net328),
    .A2(net264),
    .B1(net230),
    .B2(net1261),
    .X(_0418_));
 sky130_fd_sc_hd__a22o_1 _5315_ (.A1(net323),
    .A2(net264),
    .B1(net230),
    .B2(net1111),
    .X(_0419_));
 sky130_fd_sc_hd__a22o_1 _5316_ (.A1(net325),
    .A2(net264),
    .B1(net230),
    .B2(net1131),
    .X(_0420_));
 sky130_fd_sc_hd__a22o_1 _5317_ (.A1(net324),
    .A2(net264),
    .B1(net230),
    .B2(net1345),
    .X(_0421_));
 sky130_fd_sc_hd__a22o_1 _5318_ (.A1(net322),
    .A2(net263),
    .B1(net229),
    .B2(net1175),
    .X(_0422_));
 sky130_fd_sc_hd__a22o_1 _5319_ (.A1(net319),
    .A2(net264),
    .B1(net230),
    .B2(net1013),
    .X(_0423_));
 sky130_fd_sc_hd__a22o_1 _5320_ (.A1(net321),
    .A2(net263),
    .B1(net229),
    .B2(net1618),
    .X(_0424_));
 sky130_fd_sc_hd__a22o_1 _5321_ (.A1(net320),
    .A2(net263),
    .B1(net229),
    .B2(net1327),
    .X(_0425_));
 sky130_fd_sc_hd__a22o_1 _5322_ (.A1(net318),
    .A2(net264),
    .B1(net230),
    .B2(net1159),
    .X(_0426_));
 sky130_fd_sc_hd__a22o_1 _5323_ (.A1(net342),
    .A2(net263),
    .B1(net229),
    .B2(net999),
    .X(_0427_));
 sky130_fd_sc_hd__a22o_1 _5324_ (.A1(_1382_),
    .A2(net263),
    .B1(net229),
    .B2(net1105),
    .X(_0428_));
 sky130_fd_sc_hd__a22o_1 _5325_ (.A1(net341),
    .A2(net264),
    .B1(net230),
    .B2(net1399),
    .X(_0429_));
 sky130_fd_sc_hd__a22o_1 _5326_ (.A1(net343),
    .A2(net263),
    .B1(net229),
    .B2(net1283),
    .X(_0430_));
 sky130_fd_sc_hd__a22o_1 _5327_ (.A1(net338),
    .A2(net263),
    .B1(net229),
    .B2(net1466),
    .X(_0431_));
 sky130_fd_sc_hd__a22o_1 _5328_ (.A1(net340),
    .A2(net263),
    .B1(net229),
    .B2(net1367),
    .X(_0432_));
 sky130_fd_sc_hd__a22o_1 _5329_ (.A1(net339),
    .A2(net263),
    .B1(net229),
    .B2(net1043),
    .X(_0433_));
 sky130_fd_sc_hd__a22o_1 _5330_ (.A1(net337),
    .A2(net263),
    .B1(net229),
    .B2(net1411),
    .X(_0434_));
 sky130_fd_sc_hd__a22o_1 _5331_ (.A1(net334),
    .A2(net264),
    .B1(net230),
    .B2(net1319),
    .X(_0435_));
 sky130_fd_sc_hd__a22o_1 _5332_ (.A1(net336),
    .A2(net263),
    .B1(net229),
    .B2(net1668),
    .X(_0436_));
 sky130_fd_sc_hd__a22o_1 _5333_ (.A1(net335),
    .A2(net263),
    .B1(net229),
    .B2(net1526),
    .X(_0437_));
 sky130_fd_sc_hd__a22o_1 _5334_ (.A1(net333),
    .A2(net263),
    .B1(net229),
    .B2(net1279),
    .X(_0438_));
 sky130_fd_sc_hd__a22o_1 _5335_ (.A1(net346),
    .A2(net263),
    .B1(net229),
    .B2(net952),
    .X(_0439_));
 sky130_fd_sc_hd__a22o_1 _5336_ (.A1(net344),
    .A2(net263),
    .B1(net229),
    .B2(net1177),
    .X(_0440_));
 sky130_fd_sc_hd__a22o_1 _5337_ (.A1(net345),
    .A2(net264),
    .B1(net230),
    .B2(net1373),
    .X(_0441_));
 sky130_fd_sc_hd__a22o_1 _5338_ (.A1(net368),
    .A2(net263),
    .B1(net229),
    .B2(net1291),
    .X(_0442_));
 sky130_fd_sc_hd__nand2_4 _5339_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .Y(_2637_));
 sky130_fd_sc_hd__nor2_2 _5340_ (.A(_2617_),
    .B(_2637_),
    .Y(_2638_));
 sky130_fd_sc_hd__or2_2 _5341_ (.A(_2617_),
    .B(_2637_),
    .X(_2639_));
 sky130_fd_sc_hd__nor2_1 _5342_ (.A(net472),
    .B(net262),
    .Y(_2640_));
 sky130_fd_sc_hd__nand2_1 _5343_ (.A(net460),
    .B(_2639_),
    .Y(_2641_));
 sky130_fd_sc_hd__o22a_1 _5344_ (.A1(net329),
    .A2(_2639_),
    .B1(_2641_),
    .B2(net852),
    .X(_0443_));
 sky130_fd_sc_hd__o22a_1 _5345_ (.A1(net330),
    .A2(_2639_),
    .B1(_2641_),
    .B2(net1774),
    .X(_0444_));
 sky130_fd_sc_hd__o22a_1 _5346_ (.A1(net331),
    .A2(_2639_),
    .B1(_2641_),
    .B2(net1097),
    .X(_0445_));
 sky130_fd_sc_hd__o22a_1 _5347_ (.A1(net332),
    .A2(_2639_),
    .B1(_2641_),
    .B2(net954),
    .X(_0446_));
 sky130_fd_sc_hd__a22o_1 _5348_ (.A1(net327),
    .A2(net262),
    .B1(net228),
    .B2(net1155),
    .X(_0447_));
 sky130_fd_sc_hd__a22o_1 _5349_ (.A1(_1608_),
    .A2(net262),
    .B1(net228),
    .B2(net1584),
    .X(_0448_));
 sky130_fd_sc_hd__a22o_1 _5350_ (.A1(net326),
    .A2(net262),
    .B1(net228),
    .B2(net1323),
    .X(_0449_));
 sky130_fd_sc_hd__a22o_1 _5351_ (.A1(net328),
    .A2(net262),
    .B1(net228),
    .B2(net1257),
    .X(_0450_));
 sky130_fd_sc_hd__a22o_1 _5352_ (.A1(net323),
    .A2(net262),
    .B1(net228),
    .B2(net950),
    .X(_0451_));
 sky130_fd_sc_hd__a22o_1 _5353_ (.A1(net325),
    .A2(net262),
    .B1(net228),
    .B2(net1337),
    .X(_0452_));
 sky130_fd_sc_hd__a22o_1 _5354_ (.A1(net324),
    .A2(net262),
    .B1(net228),
    .B2(net1247),
    .X(_0453_));
 sky130_fd_sc_hd__a22o_1 _5355_ (.A1(net322),
    .A2(net261),
    .B1(net227),
    .B2(net1195),
    .X(_0454_));
 sky130_fd_sc_hd__a22o_1 _5356_ (.A1(net319),
    .A2(net262),
    .B1(net228),
    .B2(net923),
    .X(_0455_));
 sky130_fd_sc_hd__a22o_1 _5357_ (.A1(net321),
    .A2(net261),
    .B1(net227),
    .B2(net1518),
    .X(_0456_));
 sky130_fd_sc_hd__a22o_1 _5358_ (.A1(net320),
    .A2(net261),
    .B1(net227),
    .B2(net1355),
    .X(_0457_));
 sky130_fd_sc_hd__a22o_1 _5359_ (.A1(net318),
    .A2(net262),
    .B1(net228),
    .B2(net1049),
    .X(_0458_));
 sky130_fd_sc_hd__a22o_1 _5360_ (.A1(net342),
    .A2(net261),
    .B1(net227),
    .B2(net1223),
    .X(_0459_));
 sky130_fd_sc_hd__a22o_1 _5361_ (.A1(_1382_),
    .A2(net261),
    .B1(net227),
    .B2(net1001),
    .X(_0460_));
 sky130_fd_sc_hd__a22o_1 _5362_ (.A1(net341),
    .A2(net262),
    .B1(net228),
    .B2(net1409),
    .X(_0461_));
 sky130_fd_sc_hd__a22o_1 _5363_ (.A1(net343),
    .A2(net261),
    .B1(net227),
    .B2(net1474),
    .X(_0462_));
 sky130_fd_sc_hd__a22o_1 _5364_ (.A1(net338),
    .A2(net261),
    .B1(net227),
    .B2(net1407),
    .X(_0463_));
 sky130_fd_sc_hd__a22o_1 _5365_ (.A1(net340),
    .A2(net261),
    .B1(net227),
    .B2(net1063),
    .X(_0464_));
 sky130_fd_sc_hd__a22o_1 _5366_ (.A1(net339),
    .A2(net261),
    .B1(net227),
    .B2(net1494),
    .X(_0465_));
 sky130_fd_sc_hd__a22o_1 _5367_ (.A1(net337),
    .A2(net261),
    .B1(net227),
    .B2(net1307),
    .X(_0466_));
 sky130_fd_sc_hd__a22o_1 _5368_ (.A1(net334),
    .A2(net262),
    .B1(net228),
    .B2(net1418),
    .X(_0467_));
 sky130_fd_sc_hd__a22o_1 _5369_ (.A1(net336),
    .A2(net261),
    .B1(net227),
    .B2(net1299),
    .X(_0468_));
 sky130_fd_sc_hd__a22o_1 _5370_ (.A1(net335),
    .A2(net261),
    .B1(net227),
    .B2(net1391),
    .X(_0469_));
 sky130_fd_sc_hd__a22o_1 _5371_ (.A1(net333),
    .A2(net261),
    .B1(net227),
    .B2(net1718),
    .X(_0470_));
 sky130_fd_sc_hd__a22o_1 _5372_ (.A1(net346),
    .A2(net261),
    .B1(net227),
    .B2(net1253),
    .X(_0471_));
 sky130_fd_sc_hd__a22o_1 _5373_ (.A1(net344),
    .A2(net261),
    .B1(net227),
    .B2(net1448),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _5374_ (.A1(net345),
    .A2(net262),
    .B1(net228),
    .B2(net1674),
    .X(_0473_));
 sky130_fd_sc_hd__a22o_1 _5375_ (.A1(net368),
    .A2(net261),
    .B1(net227),
    .B2(net1083),
    .X(_0474_));
 sky130_fd_sc_hd__nor2_2 _5376_ (.A(_2613_),
    .B(_2617_),
    .Y(_2642_));
 sky130_fd_sc_hd__inv_2 _5377_ (.A(net259),
    .Y(_2643_));
 sky130_fd_sc_hd__nor2_2 _5378_ (.A(net471),
    .B(net259),
    .Y(_2644_));
 sky130_fd_sc_hd__or2_1 _5379_ (.A(net472),
    .B(net259),
    .X(_2645_));
 sky130_fd_sc_hd__a22o_1 _5380_ (.A1(net329),
    .A2(_2642_),
    .B1(net226),
    .B2(net1728),
    .X(_0475_));
 sky130_fd_sc_hd__a22o_1 _5381_ (.A1(net330),
    .A2(_2642_),
    .B1(net226),
    .B2(net1670),
    .X(_0476_));
 sky130_fd_sc_hd__o22a_1 _5382_ (.A1(net331),
    .A2(_2643_),
    .B1(_2645_),
    .B2(net790),
    .X(_0477_));
 sky130_fd_sc_hd__o22a_1 _5383_ (.A1(net332),
    .A2(_2643_),
    .B1(_2645_),
    .B2(net1933),
    .X(_0478_));
 sky130_fd_sc_hd__a22o_1 _5384_ (.A1(net327),
    .A2(net259),
    .B1(net226),
    .B2(net1069),
    .X(_0479_));
 sky130_fd_sc_hd__a22o_1 _5385_ (.A1(_1608_),
    .A2(net259),
    .B1(net226),
    .B2(net1395),
    .X(_0480_));
 sky130_fd_sc_hd__a22o_1 _5386_ (.A1(net326),
    .A2(net259),
    .B1(net226),
    .B2(net1542),
    .X(_0481_));
 sky130_fd_sc_hd__a22o_1 _5387_ (.A1(net328),
    .A2(net259),
    .B1(net226),
    .B2(net1550),
    .X(_0482_));
 sky130_fd_sc_hd__a22o_1 _5388_ (.A1(net323),
    .A2(net259),
    .B1(net226),
    .B2(net1229),
    .X(_0483_));
 sky130_fd_sc_hd__a22o_1 _5389_ (.A1(net325),
    .A2(net259),
    .B1(net226),
    .B2(net1349),
    .X(_0484_));
 sky130_fd_sc_hd__a22o_1 _5390_ (.A1(net324),
    .A2(net259),
    .B1(net226),
    .B2(net1233),
    .X(_0485_));
 sky130_fd_sc_hd__a22o_1 _5391_ (.A1(net322),
    .A2(net260),
    .B1(net225),
    .B2(net1634),
    .X(_0486_));
 sky130_fd_sc_hd__a22o_1 _5392_ (.A1(net319),
    .A2(net259),
    .B1(net226),
    .B2(net1432),
    .X(_0487_));
 sky130_fd_sc_hd__a22o_1 _5393_ (.A1(net321),
    .A2(net260),
    .B1(net225),
    .B2(net1652),
    .X(_0488_));
 sky130_fd_sc_hd__a22o_1 _5394_ (.A1(net320),
    .A2(net259),
    .B1(net225),
    .B2(net1804),
    .X(_0489_));
 sky130_fd_sc_hd__a22o_1 _5395_ (.A1(net318),
    .A2(net259),
    .B1(net226),
    .B2(net1570),
    .X(_0490_));
 sky130_fd_sc_hd__a22o_1 _5396_ (.A1(net342),
    .A2(net260),
    .B1(net225),
    .B2(net1255),
    .X(_0491_));
 sky130_fd_sc_hd__a22o_1 _5397_ (.A1(_1382_),
    .A2(net260),
    .B1(net225),
    .B2(net1694),
    .X(_0492_));
 sky130_fd_sc_hd__a22o_1 _5398_ (.A1(net341),
    .A2(net259),
    .B1(net226),
    .B2(net1690),
    .X(_0493_));
 sky130_fd_sc_hd__a22o_1 _5399_ (.A1(net343),
    .A2(net260),
    .B1(net225),
    .B2(net1171),
    .X(_0494_));
 sky130_fd_sc_hd__a22o_1 _5400_ (.A1(net338),
    .A2(net260),
    .B1(net225),
    .B2(net1468),
    .X(_0495_));
 sky130_fd_sc_hd__a22o_1 _5401_ (.A1(net340),
    .A2(net260),
    .B1(net225),
    .B2(net1632),
    .X(_0496_));
 sky130_fd_sc_hd__a22o_1 _5402_ (.A1(net339),
    .A2(net260),
    .B1(net225),
    .B2(net1534),
    .X(_0497_));
 sky130_fd_sc_hd__a22o_1 _5403_ (.A1(net337),
    .A2(net260),
    .B1(net225),
    .B2(net1624),
    .X(_0498_));
 sky130_fd_sc_hd__a22o_1 _5404_ (.A1(net334),
    .A2(net259),
    .B1(net226),
    .B2(net1325),
    .X(_0499_));
 sky130_fd_sc_hd__a22o_1 _5405_ (.A1(net336),
    .A2(net260),
    .B1(net225),
    .B2(net1578),
    .X(_0500_));
 sky130_fd_sc_hd__a22o_1 _5406_ (.A1(net335),
    .A2(net260),
    .B1(net225),
    .B2(net1640),
    .X(_0501_));
 sky130_fd_sc_hd__a22o_1 _5407_ (.A1(net333),
    .A2(net260),
    .B1(net225),
    .B2(net1249),
    .X(_0502_));
 sky130_fd_sc_hd__a22o_1 _5408_ (.A1(net346),
    .A2(net260),
    .B1(net225),
    .B2(net1644),
    .X(_0503_));
 sky130_fd_sc_hd__a22o_1 _5409_ (.A1(net344),
    .A2(net260),
    .B1(net225),
    .B2(net1814),
    .X(_0504_));
 sky130_fd_sc_hd__a22o_1 _5410_ (.A1(net345),
    .A2(net259),
    .B1(net226),
    .B2(net1610),
    .X(_0505_));
 sky130_fd_sc_hd__a22o_1 _5411_ (.A1(net368),
    .A2(net260),
    .B1(net225),
    .B2(net1329),
    .X(_0506_));
 sky130_fd_sc_hd__and2_4 _5412_ (.A(net174),
    .B(net277),
    .X(_2646_));
 sky130_fd_sc_hd__nand2_1 _5413_ (.A(net175),
    .B(net277),
    .Y(_2647_));
 sky130_fd_sc_hd__o31ai_1 _5414_ (.A1(net2124),
    .A2(net2071),
    .A3(_2137_),
    .B1(net2072),
    .Y(_2648_));
 sky130_fd_sc_hd__or3b_1 _5415_ (.A(_2137_),
    .B(net2124),
    .C_N(net2071),
    .X(_2649_));
 sky130_fd_sc_hd__nor2_1 _5416_ (.A(net2144),
    .B(_2649_),
    .Y(_2650_));
 sky130_fd_sc_hd__nor2_1 _5417_ (.A(net2048),
    .B(_2133_),
    .Y(_2651_));
 sky130_fd_sc_hd__nor2_1 _5418_ (.A(net2144),
    .B(net2071),
    .Y(_2652_));
 sky130_fd_sc_hd__a41o_1 _5419_ (.A1(_1277_),
    .A2(net2048),
    .A3(net2000),
    .A4(_2652_),
    .B1(_2650_),
    .X(_2653_));
 sky130_fd_sc_hd__o31a_1 _5420_ (.A1(_2648_),
    .A2(_2651_),
    .A3(_2653_),
    .B1(_2646_),
    .X(_0507_));
 sky130_fd_sc_hd__nor3_1 _5421_ (.A(net1990),
    .B(net1998),
    .C(net1698),
    .Y(_2654_));
 sky130_fd_sc_hd__a21oi_2 _5422_ (.A1(net2144),
    .A2(_2654_),
    .B1(_2649_),
    .Y(_2655_));
 sky130_fd_sc_hd__and2b_1 _5423_ (.A_N(net1990),
    .B(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__xor2_1 _5424_ (.A(net1998),
    .B(net1698),
    .X(_2657_));
 sky130_fd_sc_hd__nand2_1 _5425_ (.A(_2656_),
    .B(_2657_),
    .Y(_2658_));
 sky130_fd_sc_hd__nor2_4 _5426_ (.A(_2131_),
    .B(_2137_),
    .Y(_2659_));
 sky130_fd_sc_hd__and2_2 _5427_ (.A(net2124),
    .B(_2659_),
    .X(_2660_));
 sky130_fd_sc_hd__nand2_1 _5428_ (.A(net2124),
    .B(_2659_),
    .Y(_2661_));
 sky130_fd_sc_hd__and2_1 _5429_ (.A(net2144),
    .B(_2134_),
    .X(_2662_));
 sky130_fd_sc_hd__nand2_1 _5430_ (.A(net2144),
    .B(_2134_),
    .Y(_2663_));
 sky130_fd_sc_hd__or4b_1 _5431_ (.A(_2655_),
    .B(_2660_),
    .C(_2662_),
    .D_N(_3623_),
    .X(_2664_));
 sky130_fd_sc_hd__a21bo_1 _5432_ (.A1(_2650_),
    .A2(_2654_),
    .B1_N(_2664_),
    .X(_2665_));
 sky130_fd_sc_hd__nand2b_1 _5433_ (.A_N(_2665_),
    .B(_2658_),
    .Y(_2666_));
 sky130_fd_sc_hd__inv_2 _5434_ (.A(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__and2_1 _5435_ (.A(net1990),
    .B(_2655_),
    .X(_2668_));
 sky130_fd_sc_hd__nand2_1 _5436_ (.A(net1990),
    .B(_2655_),
    .Y(_2669_));
 sky130_fd_sc_hd__nand2_1 _5437_ (.A(net1998),
    .B(_2668_),
    .Y(_2670_));
 sky130_fd_sc_hd__nor3_1 _5438_ (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .B(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .C(_2661_),
    .Y(_2671_));
 sky130_fd_sc_hd__or3b_1 _5439_ (.A(_2669_),
    .B(net2197),
    .C_N(net1698),
    .X(_2672_));
 sky130_fd_sc_hd__o311a_1 _5440_ (.A1(net1990),
    .A2(net1998),
    .A3(_2661_),
    .B1(_2670_),
    .C1(_2672_),
    .X(_2673_));
 sky130_fd_sc_hd__nand3_1 _5441_ (.A(net1998),
    .B(net1698),
    .C(_2656_),
    .Y(_2674_));
 sky130_fd_sc_hd__o31a_1 _5442_ (.A1(net1998),
    .A2(net1698),
    .A3(_2669_),
    .B1(_2674_),
    .X(_2675_));
 sky130_fd_sc_hd__and3_1 _5443_ (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .B(net2202),
    .C(_2659_),
    .X(_2676_));
 sky130_fd_sc_hd__nand2_1 _5444_ (.A(net1990),
    .B(_2660_),
    .Y(_2677_));
 sky130_fd_sc_hd__o2111a_1 _5445_ (.A1(_0068_),
    .A2(_2662_),
    .B1(_2673_),
    .C1(_2675_),
    .D1(_2677_),
    .X(_2678_));
 sky130_fd_sc_hd__and3_1 _5446_ (.A(_2646_),
    .B(_2667_),
    .C(_2678_),
    .X(_0508_));
 sky130_fd_sc_hd__and3_1 _5447_ (.A(_1277_),
    .B(_2646_),
    .C(_2659_),
    .X(_0509_));
 sky130_fd_sc_hd__and3b_1 _5448_ (.A_N(net2144),
    .B(_2646_),
    .C(_2648_),
    .X(_0510_));
 sky130_fd_sc_hd__nand2_1 _5449_ (.A(net2048),
    .B(_2132_),
    .Y(_2679_));
 sky130_fd_sc_hd__nand2_2 _5450_ (.A(_2135_),
    .B(net2049),
    .Y(_2680_));
 sky130_fd_sc_hd__o21ai_1 _5451_ (.A1(_1277_),
    .A2(net2144),
    .B1(_2131_),
    .Y(_2681_));
 sky130_fd_sc_hd__o211a_1 _5452_ (.A1(_2137_),
    .A2(_2681_),
    .B1(_2133_),
    .C1(net2072),
    .X(_2682_));
 sky130_fd_sc_hd__nor2_1 _5453_ (.A(net162),
    .B(_2682_),
    .Y(_0511_));
 sky130_fd_sc_hd__and3_1 _5454_ (.A(net1117),
    .B(net174),
    .C(net276),
    .X(_0512_));
 sky130_fd_sc_hd__and3_1 _5455_ (.A(net894),
    .B(net179),
    .C(net281),
    .X(_0513_));
 sky130_fd_sc_hd__and3_1 _5456_ (.A(net838),
    .B(net179),
    .C(net287),
    .X(_0514_));
 sky130_fd_sc_hd__and3_1 _5457_ (.A(net886),
    .B(net176),
    .C(net281),
    .X(_0515_));
 sky130_fd_sc_hd__and3_1 _5458_ (.A(net882),
    .B(net178),
    .C(net282),
    .X(_0516_));
 sky130_fd_sc_hd__and3_1 _5459_ (.A(net930),
    .B(net179),
    .C(net288),
    .X(_0517_));
 sky130_fd_sc_hd__and3_1 _5460_ (.A(net762),
    .B(net179),
    .C(net287),
    .X(_0518_));
 sky130_fd_sc_hd__and3_1 _5461_ (.A(net919),
    .B(net180),
    .C(net288),
    .X(_0519_));
 sky130_fd_sc_hd__and3_1 _5462_ (.A(net901),
    .B(net176),
    .C(net282),
    .X(_0520_));
 sky130_fd_sc_hd__and3_1 _5463_ (.A(net832),
    .B(net175),
    .C(net279),
    .X(_0521_));
 sky130_fd_sc_hd__and3_1 _5464_ (.A(net834),
    .B(net179),
    .C(net287),
    .X(_0522_));
 sky130_fd_sc_hd__and3_1 _5465_ (.A(net807),
    .B(net175),
    .C(net279),
    .X(_0523_));
 sky130_fd_sc_hd__and3_1 _5466_ (.A(net1041),
    .B(net175),
    .C(net279),
    .X(_0524_));
 sky130_fd_sc_hd__and3_1 _5467_ (.A(net856),
    .B(net175),
    .C(net279),
    .X(_0525_));
 sky130_fd_sc_hd__and3_1 _5468_ (.A(net1029),
    .B(net178),
    .C(net284),
    .X(_0526_));
 sky130_fd_sc_hd__and3_1 _5469_ (.A(net608),
    .B(net178),
    .C(net280),
    .X(_0527_));
 sky130_fd_sc_hd__and3_1 _5470_ (.A(net1031),
    .B(net177),
    .C(net285),
    .X(_0528_));
 sky130_fd_sc_hd__and3_1 _5471_ (.A(net799),
    .B(net177),
    .C(net284),
    .X(_0529_));
 sky130_fd_sc_hd__and3_1 _5472_ (.A(net1125),
    .B(net172),
    .C(net275),
    .X(_0530_));
 sky130_fd_sc_hd__and3_1 _5473_ (.A(net871),
    .B(net172),
    .C(net274),
    .X(_0531_));
 sky130_fd_sc_hd__and3_1 _5474_ (.A(net948),
    .B(net172),
    .C(net275),
    .X(_0532_));
 sky130_fd_sc_hd__and3_1 _5475_ (.A(net915),
    .B(net172),
    .C(net274),
    .X(_0533_));
 sky130_fd_sc_hd__and3_1 _5476_ (.A(net820),
    .B(net172),
    .C(net275),
    .X(_0534_));
 sky130_fd_sc_hd__and3_1 _5477_ (.A(net774),
    .B(net173),
    .C(net273),
    .X(_0535_));
 sky130_fd_sc_hd__and3_1 _5478_ (.A(net764),
    .B(net171),
    .C(net273),
    .X(_0536_));
 sky130_fd_sc_hd__and3_1 _5479_ (.A(net803),
    .B(net173),
    .C(net273),
    .X(_0537_));
 sky130_fd_sc_hd__and3_1 _5480_ (.A(net983),
    .B(net171),
    .C(net276),
    .X(_0538_));
 sky130_fd_sc_hd__and3_1 _5481_ (.A(net658),
    .B(net171),
    .C(net271),
    .X(_0539_));
 sky130_fd_sc_hd__and3_1 _5482_ (.A(net1281),
    .B(net171),
    .C(net271),
    .X(_0540_));
 sky130_fd_sc_hd__and3_1 _5483_ (.A(net772),
    .B(net171),
    .C(net272),
    .X(_0541_));
 sky130_fd_sc_hd__and3_1 _5484_ (.A(net554),
    .B(net174),
    .C(net276),
    .X(_0542_));
 sky130_fd_sc_hd__and3_1 _5485_ (.A(net1135),
    .B(net182),
    .C(net283),
    .X(_0543_));
 sky130_fd_sc_hd__and3_1 _5486_ (.A(net969),
    .B(net179),
    .C(net282),
    .X(_0544_));
 sky130_fd_sc_hd__and3_1 _5487_ (.A(net725),
    .B(net176),
    .C(net282),
    .X(_0545_));
 sky130_fd_sc_hd__and3_1 _5488_ (.A(net842),
    .B(net176),
    .C(net282),
    .X(_0546_));
 sky130_fd_sc_hd__and3_1 _5489_ (.A(net840),
    .B(net176),
    .C(net282),
    .X(_0547_));
 sky130_fd_sc_hd__and3_1 _5490_ (.A(net741),
    .B(net179),
    .C(net281),
    .X(_0548_));
 sky130_fd_sc_hd__and3_1 _5491_ (.A(net788),
    .B(net180),
    .C(net287),
    .X(_0549_));
 sky130_fd_sc_hd__and3_1 _5492_ (.A(net552),
    .B(net175),
    .C(net279),
    .X(_0550_));
 sky130_fd_sc_hd__and3_1 _5493_ (.A(net822),
    .B(net176),
    .C(net279),
    .X(_0551_));
 sky130_fd_sc_hd__and3_1 _5494_ (.A(net580),
    .B(net180),
    .C(net289),
    .X(_0552_));
 sky130_fd_sc_hd__and3_1 _5495_ (.A(net878),
    .B(net177),
    .C(net284),
    .X(_0553_));
 sky130_fd_sc_hd__and3_1 _5496_ (.A(net884),
    .B(net178),
    .C(net280),
    .X(_0554_));
 sky130_fd_sc_hd__and3_1 _5497_ (.A(net792),
    .B(net180),
    .C(net288),
    .X(_0555_));
 sky130_fd_sc_hd__and3_1 _5498_ (.A(net548),
    .B(net176),
    .C(net283),
    .X(_0556_));
 sky130_fd_sc_hd__and3_1 _5499_ (.A(net1227),
    .B(net177),
    .C(net284),
    .X(_0557_));
 sky130_fd_sc_hd__and3_1 _5500_ (.A(net1077),
    .B(net180),
    .C(net288),
    .X(_0558_));
 sky130_fd_sc_hd__and3_1 _5501_ (.A(net1095),
    .B(net177),
    .C(net284),
    .X(_0559_));
 sky130_fd_sc_hd__and3_1 _5502_ (.A(net848),
    .B(net171),
    .C(net271),
    .X(_0560_));
 sky130_fd_sc_hd__and3_1 _5503_ (.A(net1061),
    .B(net183),
    .C(net275),
    .X(_0561_));
 sky130_fd_sc_hd__and3_1 _5504_ (.A(net1017),
    .B(net172),
    .C(net274),
    .X(_0562_));
 sky130_fd_sc_hd__and3_1 _5505_ (.A(net909),
    .B(net173),
    .C(net271),
    .X(_0563_));
 sky130_fd_sc_hd__and3_1 _5506_ (.A(net960),
    .B(net173),
    .C(net274),
    .X(_0564_));
 sky130_fd_sc_hd__and3_1 _5507_ (.A(net956),
    .B(net171),
    .C(net272),
    .X(_0565_));
 sky130_fd_sc_hd__and3_1 _5508_ (.A(net1085),
    .B(net172),
    .C(net274),
    .X(_0566_));
 sky130_fd_sc_hd__and3_1 _5509_ (.A(net648),
    .B(net171),
    .C(net272),
    .X(_0567_));
 sky130_fd_sc_hd__and3_1 _5510_ (.A(net875),
    .B(net171),
    .C(net271),
    .X(_0568_));
 sky130_fd_sc_hd__and3_1 _5511_ (.A(net1065),
    .B(net171),
    .C(net271),
    .X(_0569_));
 sky130_fd_sc_hd__and3_1 _5512_ (.A(net814),
    .B(net171),
    .C(net272),
    .X(_0570_));
 sky130_fd_sc_hd__and3_1 _5513_ (.A(net863),
    .B(net173),
    .C(net272),
    .X(_0571_));
 sky130_fd_sc_hd__and3_1 _5514_ (.A(net401),
    .B(net181),
    .C(net290),
    .X(_0572_));
 sky130_fd_sc_hd__and3_1 _5515_ (.A(net390),
    .B(net181),
    .C(net290),
    .X(_0573_));
 sky130_fd_sc_hd__and3_1 _5516_ (.A(net383),
    .B(net181),
    .C(net290),
    .X(_0574_));
 sky130_fd_sc_hd__and3_1 _5517_ (.A(net379),
    .B(net181),
    .C(net290),
    .X(_0575_));
 sky130_fd_sc_hd__and3_1 _5518_ (.A(net430),
    .B(net181),
    .C(net286),
    .X(_0576_));
 sky130_fd_sc_hd__and3_1 _5519_ (.A(net421),
    .B(net181),
    .C(net285),
    .X(_0577_));
 sky130_fd_sc_hd__and3_1 _5520_ (.A(net411),
    .B(net181),
    .C(net285),
    .X(_0578_));
 sky130_fd_sc_hd__and3_1 _5521_ (.A(net407),
    .B(net181),
    .C(net285),
    .X(_0579_));
 sky130_fd_sc_hd__and3_1 _5522_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[0] ),
    .B(net181),
    .C(net285),
    .X(_0580_));
 sky130_fd_sc_hd__and3_1 _5523_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[1] ),
    .B(net182),
    .C(net291),
    .X(_0581_));
 sky130_fd_sc_hd__and3_1 _5524_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[2] ),
    .B(net181),
    .C(net285),
    .X(_0582_));
 sky130_fd_sc_hd__and3_1 _5525_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[3] ),
    .B(net181),
    .C(net290),
    .X(_0583_));
 sky130_fd_sc_hd__and3_1 _5526_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[4] ),
    .B(net182),
    .C(net291),
    .X(_0584_));
 sky130_fd_sc_hd__and3_1 _5527_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[5] ),
    .B(net179),
    .C(net288),
    .X(_0585_));
 sky130_fd_sc_hd__and3_1 _5528_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[6] ),
    .B(net177),
    .C(net286),
    .X(_0586_));
 sky130_fd_sc_hd__and3_1 _5529_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[7] ),
    .B(net178),
    .C(net285),
    .X(_0587_));
 sky130_fd_sc_hd__and3_1 _5530_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[8] ),
    .B(net182),
    .C(net288),
    .X(_0588_));
 sky130_fd_sc_hd__and3_1 _5531_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[9] ),
    .B(net180),
    .C(net289),
    .X(_0589_));
 sky130_fd_sc_hd__and3_1 _5532_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[10] ),
    .B(net181),
    .C(net285),
    .X(_0590_));
 sky130_fd_sc_hd__and3_1 _5533_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[11] ),
    .B(net2085),
    .C(net277),
    .X(_0591_));
 sky130_fd_sc_hd__and3_1 _5534_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[12] ),
    .B(net180),
    .C(net289),
    .X(_0592_));
 sky130_fd_sc_hd__and3_1 _5535_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[13] ),
    .B(net177),
    .C(net286),
    .X(_0593_));
 sky130_fd_sc_hd__and3_1 _5536_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[14] ),
    .B(net178),
    .C(net283),
    .X(_0594_));
 sky130_fd_sc_hd__and3_1 _5537_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[15] ),
    .B(net180),
    .C(net288),
    .X(_0595_));
 sky130_fd_sc_hd__and3_1 _5538_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[16] ),
    .B(net177),
    .C(net284),
    .X(_0596_));
 sky130_fd_sc_hd__and3_1 _5539_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[17] ),
    .B(net2085),
    .C(net277),
    .X(_0597_));
 sky130_fd_sc_hd__and3_1 _5540_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[18] ),
    .B(net181),
    .C(net290),
    .X(_0598_));
 sky130_fd_sc_hd__and3_1 _5541_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[19] ),
    .B(net176),
    .C(net280),
    .X(_0599_));
 sky130_fd_sc_hd__and3_1 _5542_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[20] ),
    .B(net2085),
    .C(net278),
    .X(_0600_));
 sky130_fd_sc_hd__and3_1 _5543_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[21] ),
    .B(net2085),
    .C(net278),
    .X(_0601_));
 sky130_fd_sc_hd__and3_1 _5544_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[22] ),
    .B(net178),
    .C(net285),
    .X(_0602_));
 sky130_fd_sc_hd__and3_1 _5545_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[23] ),
    .B(net2085),
    .C(net278),
    .X(_0603_));
 sky130_fd_sc_hd__and3_1 _5546_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[24] ),
    .B(net182),
    .C(net290),
    .X(_0604_));
 sky130_fd_sc_hd__and3_1 _5547_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[25] ),
    .B(net2085),
    .C(net278),
    .X(_0605_));
 sky130_fd_sc_hd__and3_1 _5548_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[26] ),
    .B(net2085),
    .C(net277),
    .X(_0606_));
 sky130_fd_sc_hd__and3_1 _5549_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[27] ),
    .B(net177),
    .C(net286),
    .X(_0607_));
 sky130_fd_sc_hd__and3_1 _5550_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[28] ),
    .B(net2122),
    .C(net278),
    .X(_0608_));
 sky130_fd_sc_hd__and3_1 _5551_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[29] ),
    .B(net2122),
    .C(net278),
    .X(_0609_));
 sky130_fd_sc_hd__and3_1 _5552_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[30] ),
    .B(net182),
    .C(net290),
    .X(_0610_));
 sky130_fd_sc_hd__and3_1 _5553_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[31] ),
    .B(net177),
    .C(net277),
    .X(_0611_));
 sky130_fd_sc_hd__and3_1 _5554_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[0] ),
    .B(net181),
    .C(net290),
    .X(_0612_));
 sky130_fd_sc_hd__and3_1 _5555_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[1] ),
    .B(net182),
    .C(net291),
    .X(_0613_));
 sky130_fd_sc_hd__and3_1 _5556_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[2] ),
    .B(net181),
    .C(net286),
    .X(_0614_));
 sky130_fd_sc_hd__and3_1 _5557_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[3] ),
    .B(net182),
    .C(net290),
    .X(_0615_));
 sky130_fd_sc_hd__and3_1 _5558_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[4] ),
    .B(net180),
    .C(net289),
    .X(_0616_));
 sky130_fd_sc_hd__and3_1 _5559_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[5] ),
    .B(net180),
    .C(net288),
    .X(_0617_));
 sky130_fd_sc_hd__and3_1 _5560_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[6] ),
    .B(net178),
    .C(net285),
    .X(_0618_));
 sky130_fd_sc_hd__and3_1 _5561_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[7] ),
    .B(net177),
    .C(net285),
    .X(_0619_));
 sky130_fd_sc_hd__and3_1 _5562_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[8] ),
    .B(net179),
    .C(net283),
    .X(_0620_));
 sky130_fd_sc_hd__and3_1 _5563_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[9] ),
    .B(net180),
    .C(net289),
    .X(_0621_));
 sky130_fd_sc_hd__and3_1 _5564_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[10] ),
    .B(net182),
    .C(net288),
    .X(_0622_));
 sky130_fd_sc_hd__and3_1 _5565_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[11] ),
    .B(net176),
    .C(net283),
    .X(_0623_));
 sky130_fd_sc_hd__and3_1 _5566_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[12] ),
    .B(net180),
    .C(net289),
    .X(_0624_));
 sky130_fd_sc_hd__and3_1 _5567_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[13] ),
    .B(net177),
    .C(net286),
    .X(_0625_));
 sky130_fd_sc_hd__and3_1 _5568_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[14] ),
    .B(net178),
    .C(net280),
    .X(_0626_));
 sky130_fd_sc_hd__and3_1 _5569_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[15] ),
    .B(net180),
    .C(net288),
    .X(_0627_));
 sky130_fd_sc_hd__and3_1 _5570_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[16] ),
    .B(net177),
    .C(net284),
    .X(_0628_));
 sky130_fd_sc_hd__and3_1 _5571_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[17] ),
    .B(net2085),
    .C(net277),
    .X(_0629_));
 sky130_fd_sc_hd__and3_1 _5572_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[18] ),
    .B(net181),
    .C(net290),
    .X(_0630_));
 sky130_fd_sc_hd__and3_1 _5573_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[19] ),
    .B(net176),
    .C(net280),
    .X(_0631_));
 sky130_fd_sc_hd__and3_1 _5574_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[20] ),
    .B(net2085),
    .C(net278),
    .X(_0632_));
 sky130_fd_sc_hd__and3_1 _5575_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[21] ),
    .B(net2122),
    .C(net278),
    .X(_0633_));
 sky130_fd_sc_hd__and3_2 _5576_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[22] ),
    .B(net178),
    .C(net284),
    .X(_0634_));
 sky130_fd_sc_hd__and3_1 _5577_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[23] ),
    .B(net172),
    .C(net274),
    .X(_0635_));
 sky130_fd_sc_hd__and3_1 _5578_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[24] ),
    .B(net182),
    .C(net290),
    .X(_0636_));
 sky130_fd_sc_hd__and3_1 _5579_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[25] ),
    .B(net172),
    .C(net274),
    .X(_0637_));
 sky130_fd_sc_hd__and3_1 _5580_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[26] ),
    .B(net173),
    .C(net274),
    .X(_0638_));
 sky130_fd_sc_hd__and3_2 _5581_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[27] ),
    .B(net177),
    .C(net284),
    .X(_0639_));
 sky130_fd_sc_hd__and3_1 _5582_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[28] ),
    .B(net172),
    .C(net275),
    .X(_0640_));
 sky130_fd_sc_hd__and3_1 _5583_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[29] ),
    .B(net172),
    .C(net275),
    .X(_0641_));
 sky130_fd_sc_hd__and3_1 _5584_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[30] ),
    .B(net182),
    .C(net290),
    .X(_0642_));
 sky130_fd_sc_hd__and3_1 _5585_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[31] ),
    .B(net172),
    .C(net274),
    .X(_0643_));
 sky130_fd_sc_hd__and3_1 _5586_ (.A(net877),
    .B(net179),
    .C(net281),
    .X(_0644_));
 sky130_fd_sc_hd__and3_1 _5587_ (.A(net2151),
    .B(net175),
    .C(net280),
    .X(_0645_));
 sky130_fd_sc_hd__and3_1 _5588_ (.A(net2153),
    .B(net179),
    .C(net283),
    .X(_0646_));
 sky130_fd_sc_hd__and3_1 _5589_ (.A(net2107),
    .B(net182),
    .C(net283),
    .X(_0647_));
 sky130_fd_sc_hd__and3_1 _5590_ (.A(net175),
    .B(net277),
    .C(_2651_),
    .X(_0648_));
 sky130_fd_sc_hd__nor2_1 _5591_ (.A(net163),
    .B(_2661_),
    .Y(_0649_));
 sky130_fd_sc_hd__nor2_1 _5592_ (.A(_2133_),
    .B(net163),
    .Y(_0650_));
 sky130_fd_sc_hd__a21o_1 _5593_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ),
    .A2(net375),
    .B1(net1878),
    .X(_2683_));
 sky130_fd_sc_hd__and3_1 _5594_ (.A(net450),
    .B(_1790_),
    .C(net1879),
    .X(_0651_));
 sky130_fd_sc_hd__or2_1 _5595_ (.A(net467),
    .B(_1791_),
    .X(_2684_));
 sky130_fd_sc_hd__a21oi_1 _5596_ (.A1(net2138),
    .A2(_1790_),
    .B1(_2684_),
    .Y(_0652_));
 sky130_fd_sc_hd__and2_1 _5597_ (.A(net437),
    .B(_1801_),
    .X(_0653_));
 sky130_fd_sc_hd__and2_1 _5598_ (.A(net452),
    .B(net2157),
    .X(_0654_));
 sky130_fd_sc_hd__and2_1 _5599_ (.A(net451),
    .B(net2230),
    .X(_0655_));
 sky130_fd_sc_hd__and2_1 _5600_ (.A(net451),
    .B(_1820_),
    .X(_0656_));
 sky130_fd_sc_hd__and2_1 _5601_ (.A(net451),
    .B(net2173),
    .X(_0657_));
 sky130_fd_sc_hd__and2_1 _5602_ (.A(net457),
    .B(_1839_),
    .X(_0658_));
 sky130_fd_sc_hd__nor2_1 _5603_ (.A(net470),
    .B(net2163),
    .Y(_0659_));
 sky130_fd_sc_hd__and2_1 _5604_ (.A(net457),
    .B(_1858_),
    .X(_0660_));
 sky130_fd_sc_hd__and2_1 _5605_ (.A(net450),
    .B(_1867_),
    .X(_0661_));
 sky130_fd_sc_hd__and2_1 _5606_ (.A(net449),
    .B(net2192),
    .X(_0662_));
 sky130_fd_sc_hd__and2_1 _5607_ (.A(net457),
    .B(_1885_),
    .X(_0663_));
 sky130_fd_sc_hd__and2_1 _5608_ (.A(net449),
    .B(net2167),
    .X(_0664_));
 sky130_fd_sc_hd__nor2_1 _5609_ (.A(net468),
    .B(_1902_),
    .Y(_0665_));
 sky130_fd_sc_hd__and2_1 _5610_ (.A(net449),
    .B(net2196),
    .X(_0666_));
 sky130_fd_sc_hd__and2_1 _5611_ (.A(net453),
    .B(_1921_),
    .X(_0667_));
 sky130_fd_sc_hd__nor2_1 _5612_ (.A(net468),
    .B(net2078),
    .Y(_0668_));
 sky130_fd_sc_hd__and2_1 _5613_ (.A(net455),
    .B(_1939_),
    .X(_0669_));
 sky130_fd_sc_hd__and2_1 _5614_ (.A(net443),
    .B(_1948_),
    .X(_0670_));
 sky130_fd_sc_hd__nor2_1 _5615_ (.A(net467),
    .B(net2135),
    .Y(_0671_));
 sky130_fd_sc_hd__and2_1 _5616_ (.A(net442),
    .B(net2246),
    .X(_0672_));
 sky130_fd_sc_hd__nor2_1 _5617_ (.A(net464),
    .B(_1976_),
    .Y(_0673_));
 sky130_fd_sc_hd__and2_1 _5618_ (.A(net442),
    .B(net2184),
    .X(_0674_));
 sky130_fd_sc_hd__and2_1 _5619_ (.A(net441),
    .B(net2213),
    .X(_0675_));
 sky130_fd_sc_hd__and2_1 _5620_ (.A(net440),
    .B(_2003_),
    .X(_0676_));
 sky130_fd_sc_hd__and2_1 _5621_ (.A(net440),
    .B(_2012_),
    .X(_0677_));
 sky130_fd_sc_hd__and2_1 _5622_ (.A(net440),
    .B(_2021_),
    .X(_0678_));
 sky130_fd_sc_hd__and2_1 _5623_ (.A(net439),
    .B(_2030_),
    .X(_0679_));
 sky130_fd_sc_hd__and2_1 _5624_ (.A(net439),
    .B(net2043),
    .X(_0680_));
 sky130_fd_sc_hd__and2_1 _5625_ (.A(net439),
    .B(net2219),
    .X(_0681_));
 sky130_fd_sc_hd__and2_1 _5626_ (.A(net439),
    .B(net2249),
    .X(_0682_));
 sky130_fd_sc_hd__and2_1 _5627_ (.A(net2009),
    .B(net452),
    .X(_0683_));
 sky130_fd_sc_hd__and2_1 _5628_ (.A(net1868),
    .B(net452),
    .X(_0684_));
 sky130_fd_sc_hd__and2_1 _5629_ (.A(net660),
    .B(net455),
    .X(_0685_));
 sky130_fd_sc_hd__and2_1 _5630_ (.A(net743),
    .B(net455),
    .X(_0686_));
 sky130_fd_sc_hd__and2_1 _5631_ (.A(net437),
    .B(net546),
    .X(_0687_));
 sky130_fd_sc_hd__and2_1 _5632_ (.A(net451),
    .B(net666),
    .X(_0688_));
 sky130_fd_sc_hd__and2_1 _5633_ (.A(net451),
    .B(net582),
    .X(_0689_));
 sky130_fd_sc_hd__and2_1 _5634_ (.A(net451),
    .B(net588),
    .X(_0690_));
 sky130_fd_sc_hd__and2_1 _5635_ (.A(net451),
    .B(net600),
    .X(_0691_));
 sky130_fd_sc_hd__and2_1 _5636_ (.A(net457),
    .B(net602),
    .X(_0692_));
 sky130_fd_sc_hd__and2_1 _5637_ (.A(net457),
    .B(net713),
    .X(_0693_));
 sky130_fd_sc_hd__and2_1 _5638_ (.A(net458),
    .B(net707),
    .X(_0694_));
 sky130_fd_sc_hd__and2_1 _5639_ (.A(net449),
    .B(net679),
    .X(_0695_));
 sky130_fd_sc_hd__and2_1 _5640_ (.A(net443),
    .B(net780),
    .X(_0696_));
 sky130_fd_sc_hd__and2_1 _5641_ (.A(net457),
    .B(net731),
    .X(_0697_));
 sky130_fd_sc_hd__and2_1 _5642_ (.A(net449),
    .B(net576),
    .X(_0698_));
 sky130_fd_sc_hd__and2_1 _5643_ (.A(net449),
    .B(net677),
    .X(_0699_));
 sky130_fd_sc_hd__and2_1 _5644_ (.A(net449),
    .B(net614),
    .X(_0700_));
 sky130_fd_sc_hd__and2_1 _5645_ (.A(net453),
    .B(net695),
    .X(_0701_));
 sky130_fd_sc_hd__and2_1 _5646_ (.A(net450),
    .B(net729),
    .X(_0702_));
 sky130_fd_sc_hd__and2_1 _5647_ (.A(net455),
    .B(net697),
    .X(_0703_));
 sky130_fd_sc_hd__and2_1 _5648_ (.A(net447),
    .B(net566),
    .X(_0704_));
 sky130_fd_sc_hd__and2_1 _5649_ (.A(net441),
    .B(net556),
    .X(_0705_));
 sky130_fd_sc_hd__and2_1 _5650_ (.A(net442),
    .B(net715),
    .X(_0706_));
 sky130_fd_sc_hd__and2_1 _5651_ (.A(net441),
    .B(net717),
    .X(_0707_));
 sky130_fd_sc_hd__and2_1 _5652_ (.A(net442),
    .B(net752),
    .X(_0708_));
 sky130_fd_sc_hd__and2_1 _5653_ (.A(net439),
    .B(net691),
    .X(_0709_));
 sky130_fd_sc_hd__and2_1 _5654_ (.A(net440),
    .B(net650),
    .X(_0710_));
 sky130_fd_sc_hd__and2_1 _5655_ (.A(net440),
    .B(net636),
    .X(_0711_));
 sky130_fd_sc_hd__and2_1 _5656_ (.A(net440),
    .B(net656),
    .X(_0712_));
 sky130_fd_sc_hd__and2_1 _5657_ (.A(net437),
    .B(net737),
    .X(_0713_));
 sky130_fd_sc_hd__and2_1 _5658_ (.A(net437),
    .B(net754),
    .X(_0714_));
 sky130_fd_sc_hd__and2_1 _5659_ (.A(net439),
    .B(net756),
    .X(_0715_));
 sky130_fd_sc_hd__and2_1 _5660_ (.A(net439),
    .B(net735),
    .X(_0716_));
 sky130_fd_sc_hd__or3b_4 _5661_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .B(net2231),
    .C_N(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .X(_2685_));
 sky130_fd_sc_hd__nor2_8 _5662_ (.A(_1772_),
    .B(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__or2_4 _5663_ (.A(_1772_),
    .B(_2685_),
    .X(_2687_));
 sky130_fd_sc_hd__nor2_4 _5664_ (.A(_1771_),
    .B(_1775_),
    .Y(_2688_));
 sky130_fd_sc_hd__or2_4 _5665_ (.A(_1771_),
    .B(_1775_),
    .X(_2689_));
 sky130_fd_sc_hd__nor2_1 _5666_ (.A(_2686_),
    .B(_2688_),
    .Y(_2690_));
 sky130_fd_sc_hd__nand2_8 _5667_ (.A(_2687_),
    .B(_2689_),
    .Y(_2691_));
 sky130_fd_sc_hd__mux4_1 _5668_ (.A0(_1542_),
    .A1(_1569_),
    .A2(_1530_),
    .A3(_1558_),
    .S0(net200),
    .S1(net194),
    .X(_2692_));
 sky130_fd_sc_hd__mux4_1 _5669_ (.A0(_1591_),
    .A1(_1601_),
    .A2(_1616_),
    .A3(_1580_),
    .S0(net198),
    .S1(net194),
    .X(_2693_));
 sky130_fd_sc_hd__mux2_1 _5670_ (.A0(_2692_),
    .A1(_2693_),
    .S(net203),
    .X(_2694_));
 sky130_fd_sc_hd__mux2_1 _5671_ (.A0(_1638_),
    .A1(_1660_),
    .S(net192),
    .X(_2695_));
 sky130_fd_sc_hd__mux4_1 _5672_ (.A0(_1638_),
    .A1(_1660_),
    .A2(_1650_),
    .A3(_1629_),
    .S0(net192),
    .S1(net200),
    .X(_2696_));
 sky130_fd_sc_hd__mux2_1 _5673_ (.A0(_1697_),
    .A1(_1673_),
    .S(net192),
    .X(_2697_));
 sky130_fd_sc_hd__mux2_1 _5674_ (.A0(_1684_),
    .A1(_1707_),
    .S(net192),
    .X(_2698_));
 sky130_fd_sc_hd__mux2_1 _5675_ (.A0(_2697_),
    .A1(_2698_),
    .S(net197),
    .X(_2699_));
 sky130_fd_sc_hd__mux2_1 _5676_ (.A0(_2696_),
    .A1(_2699_),
    .S(net202),
    .X(_2700_));
 sky130_fd_sc_hd__mux2_1 _5677_ (.A0(_2694_),
    .A1(_2700_),
    .S(net209),
    .X(_2701_));
 sky130_fd_sc_hd__mux2_1 _5678_ (.A0(_1414_),
    .A1(_1391_),
    .S(net193),
    .X(_2702_));
 sky130_fd_sc_hd__mux2_1 _5679_ (.A0(_1425_),
    .A1(_1401_),
    .S(net193),
    .X(_2703_));
 sky130_fd_sc_hd__mux2_1 _5680_ (.A0(_2702_),
    .A1(_2703_),
    .S(net197),
    .X(_2704_));
 sky130_fd_sc_hd__mux2_1 _5681_ (.A0(_1458_),
    .A1(_1437_),
    .S(net192),
    .X(_2705_));
 sky130_fd_sc_hd__mux2_1 _5682_ (.A0(_1447_),
    .A1(_1468_),
    .S(net191),
    .X(_2706_));
 sky130_fd_sc_hd__mux2_1 _5683_ (.A0(_2705_),
    .A1(_2706_),
    .S(net196),
    .X(_2707_));
 sky130_fd_sc_hd__mux2_1 _5684_ (.A0(_2704_),
    .A1(_2707_),
    .S(net202),
    .X(_2708_));
 sky130_fd_sc_hd__mux2_1 _5685_ (.A0(_1505_),
    .A1(_1482_),
    .S(net191),
    .X(_2709_));
 sky130_fd_sc_hd__mux2_1 _5686_ (.A0(_1492_),
    .A1(_1516_),
    .S(net191),
    .X(_2710_));
 sky130_fd_sc_hd__mux2_1 _5687_ (.A0(_2709_),
    .A1(_2710_),
    .S(net196),
    .X(_2711_));
 sky130_fd_sc_hd__mux2_1 _5688_ (.A0(_1350_),
    .A1(_1373_),
    .S(net191),
    .X(_2712_));
 sky130_fd_sc_hd__mux2_1 _5689_ (.A0(_1360_),
    .A1(_1337_),
    .S(net191),
    .X(_2713_));
 sky130_fd_sc_hd__mux2_1 _5690_ (.A0(_2712_),
    .A1(_2713_),
    .S(net196),
    .X(_2714_));
 sky130_fd_sc_hd__mux2_1 _5691_ (.A0(_2711_),
    .A1(_2714_),
    .S(net201),
    .X(_2715_));
 sky130_fd_sc_hd__mux2_2 _5692_ (.A0(_2708_),
    .A1(_2715_),
    .S(net208),
    .X(_2716_));
 sky130_fd_sc_hd__mux2_1 _5693_ (.A0(_2701_),
    .A1(_2716_),
    .S(net185),
    .X(_2717_));
 sky130_fd_sc_hd__nand2_1 _5694_ (.A(_2691_),
    .B(_2717_),
    .Y(_2718_));
 sky130_fd_sc_hd__or3_1 _5695_ (.A(net210),
    .B(net203),
    .C(_1721_),
    .X(_2719_));
 sky130_fd_sc_hd__nor2_8 _5696_ (.A(_1771_),
    .B(_2685_),
    .Y(_2720_));
 sky130_fd_sc_hd__or2_4 _5697_ (.A(_1771_),
    .B(_2685_),
    .X(_2721_));
 sky130_fd_sc_hd__nor2_2 _5698_ (.A(net186),
    .B(_2721_),
    .Y(_2722_));
 sky130_fd_sc_hd__nand2_4 _5699_ (.A(net190),
    .B(_2720_),
    .Y(_2723_));
 sky130_fd_sc_hd__nor2_2 _5700_ (.A(net2356),
    .B(net2326),
    .Y(_2724_));
 sky130_fd_sc_hd__or2_1 _5701_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ),
    .X(_2725_));
 sky130_fd_sc_hd__nor2_2 _5702_ (.A(_2685_),
    .B(_2725_),
    .Y(_2726_));
 sky130_fd_sc_hd__and4bb_2 _5703_ (.A_N(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .B_N(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .C(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .D(_2724_),
    .X(_2727_));
 sky130_fd_sc_hd__or4_1 _5704_ (.A(_2691_),
    .B(_2720_),
    .C(net362),
    .D(net360),
    .X(_2728_));
 sky130_fd_sc_hd__nor2_8 _5705_ (.A(_1771_),
    .B(_1773_),
    .Y(_2729_));
 sky130_fd_sc_hd__or2_2 _5706_ (.A(_1771_),
    .B(_1773_),
    .X(_2730_));
 sky130_fd_sc_hd__a21oi_4 _5707_ (.A1(_1769_),
    .A2(_2724_),
    .B1(_2729_),
    .Y(_2731_));
 sky130_fd_sc_hd__a21o_2 _5708_ (.A1(_1769_),
    .A2(_2724_),
    .B1(_2729_),
    .X(_2732_));
 sky130_fd_sc_hd__nor2_1 _5709_ (.A(_1775_),
    .B(_2725_),
    .Y(_2733_));
 sky130_fd_sc_hd__or2_4 _5710_ (.A(_1775_),
    .B(_2725_),
    .X(_2734_));
 sky130_fd_sc_hd__nand2_1 _5711_ (.A(_2731_),
    .B(_2734_),
    .Y(_2735_));
 sky130_fd_sc_hd__and4b_1 _5712_ (.A_N(_2728_),
    .B(_2734_),
    .C(_2731_),
    .D(_1776_),
    .X(_2736_));
 sky130_fd_sc_hd__or4b_4 _5713_ (.A(_2728_),
    .B(net356),
    .C(net317),
    .D_N(_1776_),
    .X(_2737_));
 sky130_fd_sc_hd__a221o_1 _5714_ (.A1(net194),
    .A2(net360),
    .B1(_2735_),
    .B2(_1571_),
    .C1(net362),
    .X(_2738_));
 sky130_fd_sc_hd__a21oi_1 _5715_ (.A1(_1572_),
    .A2(_2738_),
    .B1(net223),
    .Y(_2739_));
 sky130_fd_sc_hd__o221a_1 _5716_ (.A1(_1766_),
    .A2(net2327),
    .B1(_2719_),
    .B2(_2723_),
    .C1(_2739_),
    .X(_2740_));
 sky130_fd_sc_hd__a221oi_4 _5717_ (.A1(_1571_),
    .A2(net223),
    .B1(net2328),
    .B2(_2718_),
    .C1(net467),
    .Y(_0717_));
 sky130_fd_sc_hd__mux2_1 _5718_ (.A0(_1437_),
    .A1(_1447_),
    .S(net193),
    .X(_2741_));
 sky130_fd_sc_hd__mux2_1 _5719_ (.A0(_1468_),
    .A1(_1505_),
    .S(net191),
    .X(_2742_));
 sky130_fd_sc_hd__mux2_1 _5720_ (.A0(_2741_),
    .A1(_2742_),
    .S(net197),
    .X(_2743_));
 sky130_fd_sc_hd__mux2_1 _5721_ (.A0(_1391_),
    .A1(_1425_),
    .S(net193),
    .X(_2744_));
 sky130_fd_sc_hd__mux2_1 _5722_ (.A0(_1401_),
    .A1(_1458_),
    .S(net193),
    .X(_2745_));
 sky130_fd_sc_hd__mux2_1 _5723_ (.A0(_2744_),
    .A1(_2745_),
    .S(net197),
    .X(_2746_));
 sky130_fd_sc_hd__mux2_1 _5724_ (.A0(_2743_),
    .A1(_2746_),
    .S(net205),
    .X(_2747_));
 sky130_fd_sc_hd__nor2_1 _5725_ (.A(net209),
    .B(_2747_),
    .Y(_2748_));
 sky130_fd_sc_hd__mux2_1 _5726_ (.A0(_1482_),
    .A1(_1492_),
    .S(net191),
    .X(_2749_));
 sky130_fd_sc_hd__mux2_1 _5727_ (.A0(_1516_),
    .A1(_1350_),
    .S(net191),
    .X(_2750_));
 sky130_fd_sc_hd__mux2_1 _5728_ (.A0(_2749_),
    .A1(_2750_),
    .S(net196),
    .X(_2751_));
 sky130_fd_sc_hd__nor2_1 _5729_ (.A(net201),
    .B(_2751_),
    .Y(_2752_));
 sky130_fd_sc_hd__and2b_1 _5730_ (.A_N(net191),
    .B(_1373_),
    .X(_2753_));
 sky130_fd_sc_hd__a21oi_1 _5731_ (.A1(_1360_),
    .A2(net191),
    .B1(_2753_),
    .Y(_2754_));
 sky130_fd_sc_hd__nor2_1 _5732_ (.A(net196),
    .B(_2754_),
    .Y(_2755_));
 sky130_fd_sc_hd__a21oi_1 _5733_ (.A1(_1337_),
    .A2(net196),
    .B1(_2755_),
    .Y(_2756_));
 sky130_fd_sc_hd__a21o_1 _5734_ (.A1(net201),
    .A2(_2756_),
    .B1(_2752_),
    .X(_2757_));
 sky130_fd_sc_hd__a21oi_1 _5735_ (.A1(net209),
    .A2(_2757_),
    .B1(_2748_),
    .Y(_2758_));
 sky130_fd_sc_hd__nor2_1 _5736_ (.A(_1338_),
    .B(net195),
    .Y(_2759_));
 sky130_fd_sc_hd__a21oi_2 _5737_ (.A1(net196),
    .A2(_2759_),
    .B1(_2755_),
    .Y(_2760_));
 sky130_fd_sc_hd__a21oi_4 _5738_ (.A1(net201),
    .A2(_2760_),
    .B1(_2752_),
    .Y(_2761_));
 sky130_fd_sc_hd__o21ba_1 _5739_ (.A1(net213),
    .A2(_2761_),
    .B1_N(_2748_),
    .X(_2762_));
 sky130_fd_sc_hd__a22o_1 _5740_ (.A1(_2686_),
    .A2(_2758_),
    .B1(_2762_),
    .B2(_2688_),
    .X(_2763_));
 sky130_fd_sc_hd__or3_1 _5741_ (.A(_1552_),
    .B(_1554_),
    .C(_2729_),
    .X(_2764_));
 sky130_fd_sc_hd__o21ai_1 _5742_ (.A1(_1552_),
    .A2(_1554_),
    .B1(_2729_),
    .Y(_2765_));
 sky130_fd_sc_hd__and3_1 _5743_ (.A(_1558_),
    .B(_2764_),
    .C(_2765_),
    .X(_2766_));
 sky130_fd_sc_hd__a21o_1 _5744_ (.A1(_2764_),
    .A2(_2765_),
    .B1(_1558_),
    .X(_2767_));
 sky130_fd_sc_hd__and2b_1 _5745_ (.A_N(_2766_),
    .B(_2767_),
    .X(_2768_));
 sky130_fd_sc_hd__mux2_1 _5746_ (.A0(_2729_),
    .A1(_1569_),
    .S(net195),
    .X(_2769_));
 sky130_fd_sc_hd__xor2_1 _5747_ (.A(_2768_),
    .B(_2769_),
    .X(_2770_));
 sky130_fd_sc_hd__a221o_1 _5748_ (.A1(_1560_),
    .A2(net362),
    .B1(net360),
    .B2(net198),
    .C1(net224),
    .X(_2771_));
 sky130_fd_sc_hd__mux2_1 _5749_ (.A0(_1558_),
    .A1(_1569_),
    .S(net194),
    .X(_2772_));
 sky130_fd_sc_hd__nand2_1 _5750_ (.A(net200),
    .B(_2772_),
    .Y(_2773_));
 sky130_fd_sc_hd__or2_1 _5751_ (.A(net203),
    .B(_2773_),
    .X(_2774_));
 sky130_fd_sc_hd__inv_2 _5752_ (.A(_2774_),
    .Y(_2775_));
 sky130_fd_sc_hd__or2_1 _5753_ (.A(net209),
    .B(_2774_),
    .X(_2776_));
 sky130_fd_sc_hd__a2bb2o_1 _5754_ (.A1_N(_2723_),
    .A2_N(_2776_),
    .B1(_2770_),
    .B2(net317),
    .X(_2777_));
 sky130_fd_sc_hd__a211o_1 _5755_ (.A1(net357),
    .A2(_2768_),
    .B1(_2771_),
    .C1(_2777_),
    .X(_2778_));
 sky130_fd_sc_hd__mux4_1 _5756_ (.A0(_1530_),
    .A1(_1558_),
    .A2(_1591_),
    .A3(_1542_),
    .S0(net200),
    .S1(net195),
    .X(_2779_));
 sky130_fd_sc_hd__mux4_1 _5757_ (.A0(_1580_),
    .A1(_1616_),
    .A2(_1650_),
    .A3(_1601_),
    .S0(net200),
    .S1(net195),
    .X(_2780_));
 sky130_fd_sc_hd__mux2_1 _5758_ (.A0(_2779_),
    .A1(_2780_),
    .S(net203),
    .X(_2781_));
 sky130_fd_sc_hd__mux2_1 _5759_ (.A0(_1673_),
    .A1(_1684_),
    .S(net192),
    .X(_2782_));
 sky130_fd_sc_hd__mux2_1 _5760_ (.A0(_1707_),
    .A1(_1414_),
    .S(net193),
    .X(_2783_));
 sky130_fd_sc_hd__mux2_1 _5761_ (.A0(_2782_),
    .A1(_2783_),
    .S(net197),
    .X(_2784_));
 sky130_fd_sc_hd__mux2_1 _5762_ (.A0(_1660_),
    .A1(_1697_),
    .S(net192),
    .X(_2785_));
 sky130_fd_sc_hd__mux4_1 _5763_ (.A0(_1629_),
    .A1(_1638_),
    .A2(_1660_),
    .A3(_1697_),
    .S0(net195),
    .S1(net198),
    .X(_2786_));
 sky130_fd_sc_hd__mux2_1 _5764_ (.A0(_2784_),
    .A1(_2786_),
    .S(_1539_),
    .X(_2787_));
 sky130_fd_sc_hd__mux2_1 _5765_ (.A0(_2781_),
    .A1(_2787_),
    .S(net210),
    .X(_2788_));
 sky130_fd_sc_hd__nor2_1 _5766_ (.A(net186),
    .B(_2690_),
    .Y(_2789_));
 sky130_fd_sc_hd__a221o_1 _5767_ (.A1(net187),
    .A2(_2763_),
    .B1(_2788_),
    .B2(_2789_),
    .C1(_2778_),
    .X(_2790_));
 sky130_fd_sc_hd__a21o_1 _5768_ (.A1(net198),
    .A2(_1558_),
    .B1(net221),
    .X(_2791_));
 sky130_fd_sc_hd__and3_1 _5769_ (.A(net443),
    .B(_2790_),
    .C(_2791_),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_1 _5770_ (.A0(_1542_),
    .A1(_1558_),
    .S(net195),
    .X(_2792_));
 sky130_fd_sc_hd__o21bai_2 _5771_ (.A1(net198),
    .A2(_2792_),
    .B1_N(_1720_),
    .Y(_2793_));
 sky130_fd_sc_hd__nor2_1 _5772_ (.A(net202),
    .B(_2793_),
    .Y(_2794_));
 sky130_fd_sc_hd__mux4_1 _5773_ (.A0(_1542_),
    .A1(_1591_),
    .A2(_1530_),
    .A3(_1616_),
    .S0(net198),
    .S1(net194),
    .X(_2795_));
 sky130_fd_sc_hd__mux4_1 _5774_ (.A0(_1601_),
    .A1(_1650_),
    .A2(_1580_),
    .A3(_1629_),
    .S0(net197),
    .S1(net192),
    .X(_2796_));
 sky130_fd_sc_hd__mux2_1 _5775_ (.A0(_2795_),
    .A1(_2796_),
    .S(net202),
    .X(_2797_));
 sky130_fd_sc_hd__mux2_1 _5776_ (.A0(_2695_),
    .A1(_2697_),
    .S(net197),
    .X(_2798_));
 sky130_fd_sc_hd__mux2_1 _5777_ (.A0(_2698_),
    .A1(_2702_),
    .S(net197),
    .X(_2799_));
 sky130_fd_sc_hd__mux2_1 _5778_ (.A0(_2798_),
    .A1(_2799_),
    .S(net202),
    .X(_2800_));
 sky130_fd_sc_hd__mux2_1 _5779_ (.A0(_2797_),
    .A1(_2800_),
    .S(net207),
    .X(_2801_));
 sky130_fd_sc_hd__a32o_1 _5780_ (.A1(net212),
    .A2(_2720_),
    .A3(_2794_),
    .B1(_2801_),
    .B2(_2691_),
    .X(_2802_));
 sky130_fd_sc_hd__and2_1 _5781_ (.A(net190),
    .B(_2802_),
    .X(_2803_));
 sky130_fd_sc_hd__mux2_1 _5782_ (.A0(_2710_),
    .A1(_2712_),
    .S(net196),
    .X(_2804_));
 sky130_fd_sc_hd__nor2_1 _5783_ (.A(net201),
    .B(_2804_),
    .Y(_2805_));
 sky130_fd_sc_hd__nand2_1 _5784_ (.A(net199),
    .B(_2713_),
    .Y(_2806_));
 sky130_fd_sc_hd__a21oi_1 _5785_ (.A1(net201),
    .A2(_2806_),
    .B1(_2805_),
    .Y(_2807_));
 sky130_fd_sc_hd__nor2_1 _5786_ (.A(net211),
    .B(_2807_),
    .Y(_2808_));
 sky130_fd_sc_hd__mux2_1 _5787_ (.A0(_2703_),
    .A1(_2705_),
    .S(net196),
    .X(_2809_));
 sky130_fd_sc_hd__mux2_1 _5788_ (.A0(_2706_),
    .A1(_2709_),
    .S(net196),
    .X(_2810_));
 sky130_fd_sc_hd__mux2_1 _5789_ (.A0(_2809_),
    .A1(_2810_),
    .S(net201),
    .X(_2811_));
 sky130_fd_sc_hd__nor2_1 _5790_ (.A(net207),
    .B(_2811_),
    .Y(_2812_));
 sky130_fd_sc_hd__or3_1 _5791_ (.A(_2689_),
    .B(_2808_),
    .C(_2812_),
    .X(_2813_));
 sky130_fd_sc_hd__o21ai_1 _5792_ (.A1(_1338_),
    .A2(net199),
    .B1(_2806_),
    .Y(_2814_));
 sky130_fd_sc_hd__o21ba_1 _5793_ (.A1(net204),
    .A2(_2814_),
    .B1_N(_2805_),
    .X(_2815_));
 sky130_fd_sc_hd__nor2_1 _5794_ (.A(net211),
    .B(_2815_),
    .Y(_2816_));
 sky130_fd_sc_hd__o31a_2 _5795_ (.A1(_2687_),
    .A2(_2812_),
    .A3(_2816_),
    .B1(_2813_),
    .X(_2817_));
 sky130_fd_sc_hd__o21a_1 _5796_ (.A1(_2766_),
    .A2(_2769_),
    .B1(_2767_),
    .X(_2818_));
 sky130_fd_sc_hd__nand2_1 _5797_ (.A(net206),
    .B(net359),
    .Y(_2819_));
 sky130_fd_sc_hd__nand2_1 _5798_ (.A(net203),
    .B(_2729_),
    .Y(_2820_));
 sky130_fd_sc_hd__and3_1 _5799_ (.A(_1542_),
    .B(_2819_),
    .C(_2820_),
    .X(_2821_));
 sky130_fd_sc_hd__a21o_1 _5800_ (.A1(_2819_),
    .A2(_2820_),
    .B1(_1542_),
    .X(_2822_));
 sky130_fd_sc_hd__and2b_1 _5801_ (.A_N(_2821_),
    .B(_2822_),
    .X(_2823_));
 sky130_fd_sc_hd__xnor2_1 _5802_ (.A(_2818_),
    .B(_2823_),
    .Y(_2824_));
 sky130_fd_sc_hd__a21oi_1 _5803_ (.A1(net203),
    .A2(net360),
    .B1(net362),
    .Y(_2825_));
 sky130_fd_sc_hd__o21a_1 _5804_ (.A1(_1543_),
    .A2(_2734_),
    .B1(_2825_),
    .X(_2826_));
 sky130_fd_sc_hd__o221a_1 _5805_ (.A1(_2731_),
    .A2(_2824_),
    .B1(_2826_),
    .B2(_1544_),
    .C1(net221),
    .X(_2827_));
 sky130_fd_sc_hd__o21ai_1 _5806_ (.A1(net190),
    .A2(_2817_),
    .B1(_2827_),
    .Y(_2828_));
 sky130_fd_sc_hd__o221a_1 _5807_ (.A1(_1543_),
    .A2(net221),
    .B1(_2803_),
    .B2(_2828_),
    .C1(net444),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _5808_ (.A0(_2741_),
    .A1(_2745_),
    .S(net199),
    .X(_2829_));
 sky130_fd_sc_hd__mux2_1 _5809_ (.A0(_2742_),
    .A1(_2749_),
    .S(net196),
    .X(_2830_));
 sky130_fd_sc_hd__mux2_1 _5810_ (.A0(_2829_),
    .A1(_2830_),
    .S(net201),
    .X(_2831_));
 sky130_fd_sc_hd__or2_1 _5811_ (.A(net196),
    .B(_2750_),
    .X(_2832_));
 sky130_fd_sc_hd__nand2_1 _5812_ (.A(net196),
    .B(_2754_),
    .Y(_2833_));
 sky130_fd_sc_hd__and3_1 _5813_ (.A(net204),
    .B(_2832_),
    .C(_2833_),
    .X(_2834_));
 sky130_fd_sc_hd__nor2_1 _5814_ (.A(_1338_),
    .B(net204),
    .Y(_2835_));
 sky130_fd_sc_hd__or2_1 _5815_ (.A(_2834_),
    .B(_2835_),
    .X(_2836_));
 sky130_fd_sc_hd__mux2_1 _5816_ (.A0(_2831_),
    .A1(_2836_),
    .S(net207),
    .X(_2837_));
 sky130_fd_sc_hd__a31oi_1 _5817_ (.A1(net201),
    .A2(net199),
    .A3(_2759_),
    .B1(_2834_),
    .Y(_2838_));
 sky130_fd_sc_hd__inv_2 _5818_ (.A(_2838_),
    .Y(_2839_));
 sky130_fd_sc_hd__mux2_1 _5819_ (.A0(_2831_),
    .A1(_2839_),
    .S(net207),
    .X(_2840_));
 sky130_fd_sc_hd__a22o_1 _5820_ (.A1(_2686_),
    .A2(_2837_),
    .B1(_2840_),
    .B2(_2688_),
    .X(_2841_));
 sky130_fd_sc_hd__xnor2_1 _5821_ (.A(net214),
    .B(_2729_),
    .Y(_2842_));
 sky130_fd_sc_hd__and2_1 _5822_ (.A(_1530_),
    .B(_2842_),
    .X(_2843_));
 sky130_fd_sc_hd__nand2_1 _5823_ (.A(_1530_),
    .B(_2842_),
    .Y(_2844_));
 sky130_fd_sc_hd__nor2_1 _5824_ (.A(_1530_),
    .B(_2842_),
    .Y(_2845_));
 sky130_fd_sc_hd__nor2_1 _5825_ (.A(_2843_),
    .B(_2845_),
    .Y(_2846_));
 sky130_fd_sc_hd__o21ai_1 _5826_ (.A1(_2818_),
    .A2(_2821_),
    .B1(_2822_),
    .Y(_2847_));
 sky130_fd_sc_hd__xnor2_1 _5827_ (.A(_2846_),
    .B(_2847_),
    .Y(_2848_));
 sky130_fd_sc_hd__mux2_1 _5828_ (.A0(_1530_),
    .A1(_1542_),
    .S(net194),
    .X(_2849_));
 sky130_fd_sc_hd__mux2_1 _5829_ (.A0(_2772_),
    .A1(_2849_),
    .S(net200),
    .X(_2850_));
 sky130_fd_sc_hd__and3_1 _5830_ (.A(net214),
    .B(net206),
    .C(_2850_),
    .X(_2851_));
 sky130_fd_sc_hd__a221o_1 _5831_ (.A1(_1531_),
    .A2(_2726_),
    .B1(net360),
    .B2(net209),
    .C1(net223),
    .X(_2852_));
 sky130_fd_sc_hd__a221o_1 _5832_ (.A1(net357),
    .A2(_2846_),
    .B1(_2851_),
    .B2(_2722_),
    .C1(_2852_),
    .X(_2853_));
 sky130_fd_sc_hd__mux4_1 _5833_ (.A0(_1530_),
    .A1(_1591_),
    .A2(_1616_),
    .A3(_1601_),
    .S0(net194),
    .S1(net198),
    .X(_2854_));
 sky130_fd_sc_hd__mux4_1 _5834_ (.A0(_1580_),
    .A1(_1629_),
    .A2(_1650_),
    .A3(_1638_),
    .S0(net197),
    .S1(net192),
    .X(_2855_));
 sky130_fd_sc_hd__mux2_1 _5835_ (.A0(_2854_),
    .A1(_2855_),
    .S(net203),
    .X(_2856_));
 sky130_fd_sc_hd__mux2_1 _5836_ (.A0(_2782_),
    .A1(_2785_),
    .S(net199),
    .X(_2857_));
 sky130_fd_sc_hd__mux2_1 _5837_ (.A0(_2744_),
    .A1(_2783_),
    .S(net199),
    .X(_2858_));
 sky130_fd_sc_hd__mux2_1 _5838_ (.A0(_2857_),
    .A1(_2858_),
    .S(net202),
    .X(_2859_));
 sky130_fd_sc_hd__mux2_1 _5839_ (.A0(_2856_),
    .A1(_2859_),
    .S(net209),
    .X(_2860_));
 sky130_fd_sc_hd__a221o_1 _5840_ (.A1(net317),
    .A2(_2848_),
    .B1(_2860_),
    .B2(_2789_),
    .C1(_2853_),
    .X(_2861_));
 sky130_fd_sc_hd__a21o_1 _5841_ (.A1(net187),
    .A2(_2841_),
    .B1(_2861_),
    .X(_2862_));
 sky130_fd_sc_hd__a21o_1 _5842_ (.A1(net209),
    .A2(_1530_),
    .B1(net221),
    .X(_2863_));
 sky130_fd_sc_hd__and3_1 _5843_ (.A(net444),
    .B(_2862_),
    .C(_2863_),
    .X(_0720_));
 sky130_fd_sc_hd__a21o_1 _5844_ (.A1(_2844_),
    .A2(_2847_),
    .B1(_2845_),
    .X(_2864_));
 sky130_fd_sc_hd__xnor2_1 _5845_ (.A(net190),
    .B(_2729_),
    .Y(_2865_));
 sky130_fd_sc_hd__nand2_1 _5846_ (.A(_1591_),
    .B(_2865_),
    .Y(_2866_));
 sky130_fd_sc_hd__nor2_1 _5847_ (.A(_1591_),
    .B(_2865_),
    .Y(_2867_));
 sky130_fd_sc_hd__or2_1 _5848_ (.A(_1591_),
    .B(_2865_),
    .X(_2868_));
 sky130_fd_sc_hd__nand2_1 _5849_ (.A(_2866_),
    .B(_2868_),
    .Y(_2869_));
 sky130_fd_sc_hd__and2_1 _5850_ (.A(_2864_),
    .B(_2869_),
    .X(_2870_));
 sky130_fd_sc_hd__nor2_1 _5851_ (.A(_2864_),
    .B(_2869_),
    .Y(_2871_));
 sky130_fd_sc_hd__mux2_1 _5852_ (.A0(_2707_),
    .A1(_2711_),
    .S(net201),
    .X(_2872_));
 sky130_fd_sc_hd__and2_2 _5853_ (.A(net204),
    .B(_2714_),
    .X(_2873_));
 sky130_fd_sc_hd__or3_1 _5854_ (.A(net211),
    .B(_2835_),
    .C(_2873_),
    .X(_2874_));
 sky130_fd_sc_hd__o21a_1 _5855_ (.A1(net207),
    .A2(_2872_),
    .B1(_2874_),
    .X(_2875_));
 sky130_fd_sc_hd__o311a_1 _5856_ (.A1(net211),
    .A2(_2686_),
    .A3(_2873_),
    .B1(_2875_),
    .C1(net184),
    .X(_2876_));
 sky130_fd_sc_hd__mux2_1 _5857_ (.A0(_2699_),
    .A1(_2704_),
    .S(net202),
    .X(_2877_));
 sky130_fd_sc_hd__mux2_1 _5858_ (.A0(_2693_),
    .A1(_2696_),
    .S(net202),
    .X(_2878_));
 sky130_fd_sc_hd__or2_1 _5859_ (.A(net209),
    .B(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__o211a_1 _5860_ (.A1(net213),
    .A2(_2877_),
    .B1(_2879_),
    .C1(net189),
    .X(_2880_));
 sky130_fd_sc_hd__o21ai_2 _5861_ (.A1(_2876_),
    .A2(_2880_),
    .B1(_2691_),
    .Y(_2881_));
 sky130_fd_sc_hd__mux4_1 _5862_ (.A0(_1542_),
    .A1(_1591_),
    .A2(_1558_),
    .A3(_1530_),
    .S0(net200),
    .S1(net194),
    .X(_2882_));
 sky130_fd_sc_hd__mux2_1 _5863_ (.A0(_1722_),
    .A1(_2882_),
    .S(net206),
    .X(_2883_));
 sky130_fd_sc_hd__nand2_1 _5864_ (.A(net213),
    .B(_2883_),
    .Y(_2884_));
 sky130_fd_sc_hd__inv_2 _5865_ (.A(_2884_),
    .Y(_2885_));
 sky130_fd_sc_hd__a221o_1 _5866_ (.A1(net187),
    .A2(net360),
    .B1(net357),
    .B2(_1592_),
    .C1(net362),
    .X(_2886_));
 sky130_fd_sc_hd__nand2_1 _5867_ (.A(_1593_),
    .B(_2886_),
    .Y(_2887_));
 sky130_fd_sc_hd__o211a_1 _5868_ (.A1(_2723_),
    .A2(_2884_),
    .B1(_2887_),
    .C1(net221),
    .X(_2888_));
 sky130_fd_sc_hd__o311a_1 _5869_ (.A1(_2731_),
    .A2(_2870_),
    .A3(_2871_),
    .B1(_2881_),
    .C1(_2888_),
    .X(_2889_));
 sky130_fd_sc_hd__a211oi_1 _5870_ (.A1(_1592_),
    .A2(net223),
    .B1(_2889_),
    .C1(net467),
    .Y(_0721_));
 sky130_fd_sc_hd__xnor2_1 _5871_ (.A(_1614_),
    .B(net359),
    .Y(_2890_));
 sky130_fd_sc_hd__nor2_1 _5872_ (.A(_1616_),
    .B(_2890_),
    .Y(_2891_));
 sky130_fd_sc_hd__nand2_1 _5873_ (.A(_1616_),
    .B(_2890_),
    .Y(_2892_));
 sky130_fd_sc_hd__and2b_1 _5874_ (.A_N(_2891_),
    .B(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__a21o_1 _5875_ (.A1(_2864_),
    .A2(_2866_),
    .B1(_2867_),
    .X(_2894_));
 sky130_fd_sc_hd__xnor2_1 _5876_ (.A(_2893_),
    .B(_2894_),
    .Y(_2895_));
 sky130_fd_sc_hd__mux2_1 _5877_ (.A0(_2743_),
    .A1(_2751_),
    .S(net202),
    .X(_2896_));
 sky130_fd_sc_hd__nor2_1 _5878_ (.A(net208),
    .B(_2896_),
    .Y(_2897_));
 sky130_fd_sc_hd__nor2_1 _5879_ (.A(net201),
    .B(_2760_),
    .Y(_2898_));
 sky130_fd_sc_hd__inv_2 _5880_ (.A(_2898_),
    .Y(_2899_));
 sky130_fd_sc_hd__a211o_1 _5881_ (.A1(net208),
    .A2(_2899_),
    .B1(_2897_),
    .C1(_2689_),
    .X(_2900_));
 sky130_fd_sc_hd__o21ba_1 _5882_ (.A1(net201),
    .A2(_2756_),
    .B1_N(_2835_),
    .X(_2901_));
 sky130_fd_sc_hd__a21oi_1 _5883_ (.A1(net208),
    .A2(_2901_),
    .B1(_2897_),
    .Y(_2902_));
 sky130_fd_sc_hd__nand2_1 _5884_ (.A(_2686_),
    .B(_2902_),
    .Y(_2903_));
 sky130_fd_sc_hd__a21oi_4 _5885_ (.A1(_2900_),
    .A2(_2903_),
    .B1(net189),
    .Y(_2904_));
 sky130_fd_sc_hd__a221o_1 _5886_ (.A1(_1617_),
    .A2(net362),
    .B1(net360),
    .B2(_1614_),
    .C1(net223),
    .X(_2905_));
 sky130_fd_sc_hd__a21o_1 _5887_ (.A1(net357),
    .A2(_2893_),
    .B1(_2905_),
    .X(_2906_));
 sky130_fd_sc_hd__mux2_1 _5888_ (.A0(_1616_),
    .A1(_1591_),
    .S(net194),
    .X(_2907_));
 sky130_fd_sc_hd__or2_1 _5889_ (.A(net198),
    .B(_2907_),
    .X(_2908_));
 sky130_fd_sc_hd__o21ai_1 _5890_ (.A1(net200),
    .A2(_2849_),
    .B1(_2908_),
    .Y(_2909_));
 sky130_fd_sc_hd__mux2_1 _5891_ (.A0(_2773_),
    .A1(_2909_),
    .S(net206),
    .X(_2910_));
 sky130_fd_sc_hd__mux2_1 _5892_ (.A0(_2780_),
    .A1(_2786_),
    .S(net203),
    .X(_2911_));
 sky130_fd_sc_hd__mux2_1 _5893_ (.A0(_2746_),
    .A1(_2784_),
    .S(net205),
    .X(_2912_));
 sky130_fd_sc_hd__mux2_1 _5894_ (.A0(_2911_),
    .A1(_2912_),
    .S(net210),
    .X(_2913_));
 sky130_fd_sc_hd__inv_2 _5895_ (.A(_2913_),
    .Y(_2914_));
 sky130_fd_sc_hd__o32a_1 _5896_ (.A1(net210),
    .A2(_2721_),
    .A3(_2910_),
    .B1(_2914_),
    .B2(_2690_),
    .X(_2915_));
 sky130_fd_sc_hd__a2bb2o_1 _5897_ (.A1_N(net187),
    .A2_N(_2915_),
    .B1(_2895_),
    .B2(net317),
    .X(_2916_));
 sky130_fd_sc_hd__a21oi_1 _5898_ (.A1(_1618_),
    .A2(net223),
    .B1(net467),
    .Y(_2917_));
 sky130_fd_sc_hd__o31a_2 _5899_ (.A1(_2904_),
    .A2(_2906_),
    .A3(_2916_),
    .B1(_2917_),
    .X(_0722_));
 sky130_fd_sc_hd__a21o_1 _5900_ (.A1(_2892_),
    .A2(_2894_),
    .B1(_2891_),
    .X(_2918_));
 sky130_fd_sc_hd__xnor2_1 _5901_ (.A(_1599_),
    .B(net359),
    .Y(_2919_));
 sky130_fd_sc_hd__nand2_1 _5902_ (.A(_1601_),
    .B(_2919_),
    .Y(_2920_));
 sky130_fd_sc_hd__nor2_1 _5903_ (.A(_1601_),
    .B(_2919_),
    .Y(_2921_));
 sky130_fd_sc_hd__or2_1 _5904_ (.A(_1601_),
    .B(_2919_),
    .X(_2922_));
 sky130_fd_sc_hd__nand2_1 _5905_ (.A(_2920_),
    .B(_2922_),
    .Y(_2923_));
 sky130_fd_sc_hd__a21o_1 _5906_ (.A1(_2918_),
    .A2(_2923_),
    .B1(_2731_),
    .X(_2924_));
 sky130_fd_sc_hd__o21bai_1 _5907_ (.A1(_2918_),
    .A2(_2923_),
    .B1_N(_2924_),
    .Y(_2925_));
 sky130_fd_sc_hd__a221o_1 _5908_ (.A1(_1599_),
    .A2(net360),
    .B1(net357),
    .B2(_1602_),
    .C1(net362),
    .X(_2926_));
 sky130_fd_sc_hd__o21ai_1 _5909_ (.A1(_1599_),
    .A2(_1601_),
    .B1(_2926_),
    .Y(_2927_));
 sky130_fd_sc_hd__mux2_1 _5910_ (.A0(_2796_),
    .A1(_2798_),
    .S(net202),
    .X(_2928_));
 sky130_fd_sc_hd__mux2_1 _5911_ (.A0(_2799_),
    .A1(_2809_),
    .S(net201),
    .X(_2929_));
 sky130_fd_sc_hd__mux2_1 _5912_ (.A0(_2928_),
    .A1(_2929_),
    .S(net208),
    .X(_2930_));
 sky130_fd_sc_hd__nand2_1 _5913_ (.A(_2691_),
    .B(_2930_),
    .Y(_2931_));
 sky130_fd_sc_hd__mux4_2 _5914_ (.A0(_1591_),
    .A1(_1601_),
    .A2(_1530_),
    .A3(_1616_),
    .S0(net200),
    .S1(net194),
    .X(_2932_));
 sky130_fd_sc_hd__inv_2 _5915_ (.A(_2932_),
    .Y(_2933_));
 sky130_fd_sc_hd__mux2_1 _5916_ (.A0(_2793_),
    .A1(_2933_),
    .S(net205),
    .X(_2934_));
 sky130_fd_sc_hd__or3_1 _5917_ (.A(net208),
    .B(_2721_),
    .C(_2934_),
    .X(_2935_));
 sky130_fd_sc_hd__mux2_1 _5918_ (.A0(_2804_),
    .A1(_2810_),
    .S(net204),
    .X(_2936_));
 sky130_fd_sc_hd__or2_1 _5919_ (.A(net207),
    .B(_2936_),
    .X(_2937_));
 sky130_fd_sc_hd__a21o_1 _5920_ (.A1(net204),
    .A2(_2814_),
    .B1(_2835_),
    .X(_2938_));
 sky130_fd_sc_hd__o21ai_1 _5921_ (.A1(net211),
    .A2(_2938_),
    .B1(_2937_),
    .Y(_2939_));
 sky130_fd_sc_hd__nor2_2 _5922_ (.A(net207),
    .B(_2689_),
    .Y(_2940_));
 sky130_fd_sc_hd__nand2_1 _5923_ (.A(net211),
    .B(_2688_),
    .Y(_2941_));
 sky130_fd_sc_hd__nor2_1 _5924_ (.A(net201),
    .B(_2806_),
    .Y(_2942_));
 sky130_fd_sc_hd__inv_2 _5925_ (.A(_2942_),
    .Y(_2943_));
 sky130_fd_sc_hd__o211a_1 _5926_ (.A1(net211),
    .A2(_2942_),
    .B1(_2937_),
    .C1(_2688_),
    .X(_2944_));
 sky130_fd_sc_hd__inv_2 _5927_ (.A(_2944_),
    .Y(_2945_));
 sky130_fd_sc_hd__o211a_1 _5928_ (.A1(_2687_),
    .A2(_2939_),
    .B1(_2945_),
    .C1(net184),
    .X(_2946_));
 sky130_fd_sc_hd__a31o_2 _5929_ (.A1(net189),
    .A2(_2931_),
    .A3(_2935_),
    .B1(_2946_),
    .X(_2947_));
 sky130_fd_sc_hd__and3_1 _5930_ (.A(net221),
    .B(_2927_),
    .C(_2947_),
    .X(_2948_));
 sky130_fd_sc_hd__a221oi_1 _5931_ (.A1(_1602_),
    .A2(net224),
    .B1(_2925_),
    .B2(_2948_),
    .C1(net467),
    .Y(_0723_));
 sky130_fd_sc_hd__xnor2_1 _5932_ (.A(_1578_),
    .B(net358),
    .Y(_2949_));
 sky130_fd_sc_hd__nor2_1 _5933_ (.A(_1580_),
    .B(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__nand2_1 _5934_ (.A(_1580_),
    .B(_2949_),
    .Y(_2951_));
 sky130_fd_sc_hd__nand2b_1 _5935_ (.A_N(_2950_),
    .B(_2951_),
    .Y(_2952_));
 sky130_fd_sc_hd__a21o_1 _5936_ (.A1(_2918_),
    .A2(_2920_),
    .B1(_2921_),
    .X(_2953_));
 sky130_fd_sc_hd__xnor2_1 _5937_ (.A(_2952_),
    .B(_2953_),
    .Y(_2954_));
 sky130_fd_sc_hd__nor2_1 _5938_ (.A(_2731_),
    .B(_2954_),
    .Y(_2955_));
 sky130_fd_sc_hd__mux2_1 _5939_ (.A0(_1580_),
    .A1(_1601_),
    .S(net192),
    .X(_2956_));
 sky130_fd_sc_hd__mux2_1 _5940_ (.A0(_2907_),
    .A1(_2956_),
    .S(net200),
    .X(_2957_));
 sky130_fd_sc_hd__mux2_1 _5941_ (.A0(_2850_),
    .A1(_2957_),
    .S(net205),
    .X(_2958_));
 sky130_fd_sc_hd__and3_1 _5942_ (.A(net212),
    .B(_2720_),
    .C(_2958_),
    .X(_2959_));
 sky130_fd_sc_hd__mux2_1 _5943_ (.A0(_2855_),
    .A1(_2857_),
    .S(net202),
    .X(_2960_));
 sky130_fd_sc_hd__mux2_1 _5944_ (.A0(_2829_),
    .A1(_2858_),
    .S(net204),
    .X(_2961_));
 sky130_fd_sc_hd__mux2_1 _5945_ (.A0(_2960_),
    .A1(_2961_),
    .S(net207),
    .X(_2962_));
 sky130_fd_sc_hd__a21o_1 _5946_ (.A1(_2691_),
    .A2(_2962_),
    .B1(_2959_),
    .X(_2963_));
 sky130_fd_sc_hd__o21a_1 _5947_ (.A1(_1578_),
    .A2(_1580_),
    .B1(net363),
    .X(_2964_));
 sky130_fd_sc_hd__a2bb2o_1 _5948_ (.A1_N(_2734_),
    .A2_N(_2952_),
    .B1(_2963_),
    .B2(net188),
    .X(_2965_));
 sky130_fd_sc_hd__a2111o_1 _5949_ (.A1(_1578_),
    .A2(net361),
    .B1(net222),
    .C1(_2964_),
    .D1(_2965_),
    .X(_2966_));
 sky130_fd_sc_hd__and2_1 _5950_ (.A(net204),
    .B(_2830_),
    .X(_2967_));
 sky130_fd_sc_hd__a31o_1 _5951_ (.A1(net201),
    .A2(_2832_),
    .A3(_2833_),
    .B1(_2967_),
    .X(_2968_));
 sky130_fd_sc_hd__or2_1 _5952_ (.A(net207),
    .B(_2968_),
    .X(_2969_));
 sky130_fd_sc_hd__and3_1 _5953_ (.A(net204),
    .B(net199),
    .C(_2759_),
    .X(_2970_));
 sky130_fd_sc_hd__o211a_1 _5954_ (.A1(net212),
    .A2(_2970_),
    .B1(_2969_),
    .C1(_2688_),
    .X(_2971_));
 sky130_fd_sc_hd__o21ai_1 _5955_ (.A1(_1337_),
    .A2(net211),
    .B1(_2969_),
    .Y(_2972_));
 sky130_fd_sc_hd__nor2_1 _5956_ (.A(_2687_),
    .B(_2972_),
    .Y(_2973_));
 sky130_fd_sc_hd__o21a_1 _5957_ (.A1(_2971_),
    .A2(_2973_),
    .B1(net184),
    .X(_2974_));
 sky130_fd_sc_hd__a21o_1 _5958_ (.A1(_1578_),
    .A2(_1580_),
    .B1(net221),
    .X(_2975_));
 sky130_fd_sc_hd__o311a_1 _5959_ (.A1(_2955_),
    .A2(_2966_),
    .A3(_2974_),
    .B1(_2975_),
    .C1(net438),
    .X(_0724_));
 sky130_fd_sc_hd__a21o_1 _5960_ (.A1(_2951_),
    .A2(_2953_),
    .B1(_2950_),
    .X(_2976_));
 sky130_fd_sc_hd__xnor2_1 _5961_ (.A(_1648_),
    .B(net358),
    .Y(_2977_));
 sky130_fd_sc_hd__nand2_1 _5962_ (.A(_1650_),
    .B(_2977_),
    .Y(_2978_));
 sky130_fd_sc_hd__nor2_1 _5963_ (.A(_1650_),
    .B(_2977_),
    .Y(_2979_));
 sky130_fd_sc_hd__inv_2 _5964_ (.A(_2979_),
    .Y(_2980_));
 sky130_fd_sc_hd__nand2_1 _5965_ (.A(_2978_),
    .B(_2980_),
    .Y(_2981_));
 sky130_fd_sc_hd__xor2_1 _5966_ (.A(_2976_),
    .B(_2981_),
    .X(_2982_));
 sky130_fd_sc_hd__mux4_1 _5967_ (.A0(_1601_),
    .A1(_1650_),
    .A2(_1616_),
    .A3(_1580_),
    .S0(net200),
    .S1(net194),
    .X(_2983_));
 sky130_fd_sc_hd__mux2_1 _5968_ (.A0(_2882_),
    .A1(_2983_),
    .S(net206),
    .X(_2984_));
 sky130_fd_sc_hd__o21ai_1 _5969_ (.A1(net203),
    .A2(_1721_),
    .B1(net210),
    .Y(_2985_));
 sky130_fd_sc_hd__o211ai_2 _5970_ (.A1(net209),
    .A2(_2984_),
    .B1(_2985_),
    .C1(_2720_),
    .Y(_2986_));
 sky130_fd_sc_hd__mux2_1 _5971_ (.A0(_2700_),
    .A1(_2708_),
    .S(net209),
    .X(_2987_));
 sky130_fd_sc_hd__a21bo_1 _5972_ (.A1(_2691_),
    .A2(_2987_),
    .B1_N(_2986_),
    .X(_2988_));
 sky130_fd_sc_hd__nor2_2 _5973_ (.A(_1338_),
    .B(net211),
    .Y(_2989_));
 sky130_fd_sc_hd__and2_1 _5974_ (.A(net211),
    .B(_2715_),
    .X(_2990_));
 sky130_fd_sc_hd__a22o_1 _5975_ (.A1(_2686_),
    .A2(_2989_),
    .B1(_2990_),
    .B2(_2691_),
    .X(_2991_));
 sky130_fd_sc_hd__a221o_1 _5976_ (.A1(_1648_),
    .A2(net361),
    .B1(net356),
    .B2(_1651_),
    .C1(net363),
    .X(_2992_));
 sky130_fd_sc_hd__o21a_1 _5977_ (.A1(_1648_),
    .A2(_1650_),
    .B1(_2992_),
    .X(_2993_));
 sky130_fd_sc_hd__a211o_1 _5978_ (.A1(net185),
    .A2(_2991_),
    .B1(_2993_),
    .C1(net224),
    .X(_2994_));
 sky130_fd_sc_hd__a221o_1 _5979_ (.A1(_2732_),
    .A2(_2982_),
    .B1(_2988_),
    .B2(net189),
    .C1(_2994_),
    .X(_2995_));
 sky130_fd_sc_hd__nand2_1 _5980_ (.A(_1651_),
    .B(net224),
    .Y(_2996_));
 sky130_fd_sc_hd__and3_1 _5981_ (.A(net438),
    .B(_2995_),
    .C(_2996_),
    .X(_0725_));
 sky130_fd_sc_hd__xnor2_1 _5982_ (.A(_1627_),
    .B(net358),
    .Y(_2997_));
 sky130_fd_sc_hd__and2_1 _5983_ (.A(_1629_),
    .B(_2997_),
    .X(_2998_));
 sky130_fd_sc_hd__nand2_1 _5984_ (.A(_1629_),
    .B(_2997_),
    .Y(_2999_));
 sky130_fd_sc_hd__nor2_1 _5985_ (.A(_1629_),
    .B(_2997_),
    .Y(_3000_));
 sky130_fd_sc_hd__nor2_1 _5986_ (.A(_2998_),
    .B(_3000_),
    .Y(_3001_));
 sky130_fd_sc_hd__a21o_1 _5987_ (.A1(_2976_),
    .A2(_2978_),
    .B1(_2979_),
    .X(_3002_));
 sky130_fd_sc_hd__xor2_1 _5988_ (.A(_3001_),
    .B(_3002_),
    .X(_3003_));
 sky130_fd_sc_hd__or2_1 _5989_ (.A(net206),
    .B(_2909_),
    .X(_3004_));
 sky130_fd_sc_hd__mux2_1 _5990_ (.A0(_1629_),
    .A1(_1650_),
    .S(net192),
    .X(_3005_));
 sky130_fd_sc_hd__or2_1 _5991_ (.A(net197),
    .B(_3005_),
    .X(_3006_));
 sky130_fd_sc_hd__o21ai_1 _5992_ (.A1(net200),
    .A2(_2956_),
    .B1(_3006_),
    .Y(_3007_));
 sky130_fd_sc_hd__o21ai_1 _5993_ (.A1(net203),
    .A2(_3007_),
    .B1(_3004_),
    .Y(_3008_));
 sky130_fd_sc_hd__mux2_1 _5994_ (.A0(_2775_),
    .A1(_3008_),
    .S(net214),
    .X(_3009_));
 sky130_fd_sc_hd__mux2_1 _5995_ (.A0(_2747_),
    .A1(_2787_),
    .S(net213),
    .X(_3010_));
 sky130_fd_sc_hd__a22o_1 _5996_ (.A1(_2720_),
    .A2(_3009_),
    .B1(_3010_),
    .B2(_2691_),
    .X(_3011_));
 sky130_fd_sc_hd__o21a_1 _5997_ (.A1(_1627_),
    .A2(_1629_),
    .B1(net363),
    .X(_3012_));
 sky130_fd_sc_hd__a22o_1 _5998_ (.A1(net356),
    .A2(_3001_),
    .B1(_3011_),
    .B2(net189),
    .X(_3013_));
 sky130_fd_sc_hd__a2111o_1 _5999_ (.A1(_1627_),
    .A2(net361),
    .B1(net224),
    .C1(_3012_),
    .D1(_3013_),
    .X(_3014_));
 sky130_fd_sc_hd__mux2_1 _6000_ (.A0(_1338_),
    .A1(_2757_),
    .S(net212),
    .X(_3015_));
 sky130_fd_sc_hd__o2bb2a_1 _6001_ (.A1_N(_2761_),
    .A2_N(_2940_),
    .B1(_3015_),
    .B2(_2687_),
    .X(_3016_));
 sky130_fd_sc_hd__o22ai_1 _6002_ (.A1(_2731_),
    .A2(_3003_),
    .B1(_3016_),
    .B2(net189),
    .Y(_3017_));
 sky130_fd_sc_hd__a21o_1 _6003_ (.A1(_1627_),
    .A2(_1629_),
    .B1(net221),
    .X(_3018_));
 sky130_fd_sc_hd__o211a_1 _6004_ (.A1(_3014_),
    .A2(_3017_),
    .B1(net2337),
    .C1(net438),
    .X(_0726_));
 sky130_fd_sc_hd__a21o_1 _6005_ (.A1(_2999_),
    .A2(_3002_),
    .B1(_3000_),
    .X(_3019_));
 sky130_fd_sc_hd__xnor2_1 _6006_ (.A(_1636_),
    .B(net358),
    .Y(_3020_));
 sky130_fd_sc_hd__nand2_1 _6007_ (.A(_1638_),
    .B(_3020_),
    .Y(_3021_));
 sky130_fd_sc_hd__nor2_1 _6008_ (.A(_1638_),
    .B(_3020_),
    .Y(_3022_));
 sky130_fd_sc_hd__inv_2 _6009_ (.A(_3022_),
    .Y(_3023_));
 sky130_fd_sc_hd__a21bo_1 _6010_ (.A1(_3021_),
    .A2(_3023_),
    .B1_N(_3019_),
    .X(_3024_));
 sky130_fd_sc_hd__or3b_1 _6011_ (.A(_3022_),
    .B(_3019_),
    .C_N(_3021_),
    .X(_3025_));
 sky130_fd_sc_hd__mux4_1 _6012_ (.A0(_1638_),
    .A1(_1650_),
    .A2(_1629_),
    .A3(_1580_),
    .S0(net197),
    .S1(net192),
    .X(_3026_));
 sky130_fd_sc_hd__mux2_1 _6013_ (.A0(_2932_),
    .A1(_3026_),
    .S(net205),
    .X(_3027_));
 sky130_fd_sc_hd__mux2_1 _6014_ (.A0(_2794_),
    .A1(_3027_),
    .S(net212),
    .X(_3028_));
 sky130_fd_sc_hd__nand2_1 _6015_ (.A(_2720_),
    .B(_3028_),
    .Y(_3029_));
 sky130_fd_sc_hd__mux2_1 _6016_ (.A0(_2800_),
    .A1(_2811_),
    .S(net207),
    .X(_3030_));
 sky130_fd_sc_hd__nand2_1 _6017_ (.A(_2691_),
    .B(_3030_),
    .Y(_3031_));
 sky130_fd_sc_hd__a21oi_1 _6018_ (.A1(_3029_),
    .A2(_3031_),
    .B1(net184),
    .Y(_3032_));
 sky130_fd_sc_hd__a221o_1 _6019_ (.A1(_1636_),
    .A2(net361),
    .B1(net356),
    .B2(_1639_),
    .C1(net363),
    .X(_3033_));
 sky130_fd_sc_hd__nand2_1 _6020_ (.A(_2807_),
    .B(_2940_),
    .Y(_3034_));
 sky130_fd_sc_hd__a21oi_1 _6021_ (.A1(net211),
    .A2(_2815_),
    .B1(_2989_),
    .Y(_3035_));
 sky130_fd_sc_hd__o21ai_1 _6022_ (.A1(_2687_),
    .A2(_3035_),
    .B1(_3034_),
    .Y(_3036_));
 sky130_fd_sc_hd__a221o_1 _6023_ (.A1(_1640_),
    .A2(_3033_),
    .B1(_3036_),
    .B2(net184),
    .C1(net222),
    .X(_3037_));
 sky130_fd_sc_hd__a311oi_4 _6024_ (.A1(net317),
    .A2(_3024_),
    .A3(_3025_),
    .B1(_3032_),
    .C1(_3037_),
    .Y(_3038_));
 sky130_fd_sc_hd__a211oi_4 _6025_ (.A1(_1639_),
    .A2(net224),
    .B1(_3038_),
    .C1(net466),
    .Y(_0727_));
 sky130_fd_sc_hd__xnor2_1 _6026_ (.A(_1658_),
    .B(net358),
    .Y(_3039_));
 sky130_fd_sc_hd__and2_1 _6027_ (.A(_1660_),
    .B(_3039_),
    .X(_3040_));
 sky130_fd_sc_hd__nand2_1 _6028_ (.A(_1660_),
    .B(_3039_),
    .Y(_3041_));
 sky130_fd_sc_hd__nor2_1 _6029_ (.A(_1660_),
    .B(_3039_),
    .Y(_3042_));
 sky130_fd_sc_hd__nor2_1 _6030_ (.A(_3040_),
    .B(_3042_),
    .Y(_3043_));
 sky130_fd_sc_hd__a21o_1 _6031_ (.A1(_3019_),
    .A2(_3021_),
    .B1(_3022_),
    .X(_3044_));
 sky130_fd_sc_hd__xnor2_1 _6032_ (.A(_3043_),
    .B(_3044_),
    .Y(_3045_));
 sky130_fd_sc_hd__mux4_1 _6033_ (.A0(_1629_),
    .A1(_1650_),
    .A2(_1660_),
    .A3(_1638_),
    .S0(net192),
    .S1(net199),
    .X(_3046_));
 sky130_fd_sc_hd__mux2_1 _6034_ (.A0(_2957_),
    .A1(_3046_),
    .S(net205),
    .X(_3047_));
 sky130_fd_sc_hd__a21o_1 _6035_ (.A1(net205),
    .A2(_2850_),
    .B1(net212),
    .X(_3048_));
 sky130_fd_sc_hd__o211ai_2 _6036_ (.A1(net208),
    .A2(_3047_),
    .B1(_3048_),
    .C1(_2720_),
    .Y(_3049_));
 sky130_fd_sc_hd__mux2_1 _6037_ (.A0(_2831_),
    .A1(_2859_),
    .S(net211),
    .X(_3050_));
 sky130_fd_sc_hd__a21bo_1 _6038_ (.A1(_2691_),
    .A2(_3050_),
    .B1_N(_3049_),
    .X(_3051_));
 sky130_fd_sc_hd__a221o_1 _6039_ (.A1(_1661_),
    .A2(net363),
    .B1(net361),
    .B2(_1658_),
    .C1(net222),
    .X(_3052_));
 sky130_fd_sc_hd__a22o_1 _6040_ (.A1(net356),
    .A2(_3043_),
    .B1(_3051_),
    .B2(net188),
    .X(_3053_));
 sky130_fd_sc_hd__a21oi_1 _6041_ (.A1(net212),
    .A2(_2836_),
    .B1(_2989_),
    .Y(_3054_));
 sky130_fd_sc_hd__a2bb2o_1 _6042_ (.A1_N(_2687_),
    .A2_N(_3054_),
    .B1(_2940_),
    .B2(_2839_),
    .X(_3055_));
 sky130_fd_sc_hd__a22o_1 _6043_ (.A1(net317),
    .A2(_3045_),
    .B1(_3055_),
    .B2(net184),
    .X(_3056_));
 sky130_fd_sc_hd__a21oi_1 _6044_ (.A1(_1658_),
    .A2(_1660_),
    .B1(net221),
    .Y(_3057_));
 sky130_fd_sc_hd__nor2_1 _6045_ (.A(net466),
    .B(_3057_),
    .Y(_3058_));
 sky130_fd_sc_hd__o31a_1 _6046_ (.A1(_3052_),
    .A2(_3053_),
    .A3(_3056_),
    .B1(_3058_),
    .X(_0728_));
 sky130_fd_sc_hd__a21o_2 _6047_ (.A1(_3041_),
    .A2(_3044_),
    .B1(_3042_),
    .X(_3059_));
 sky130_fd_sc_hd__xnor2_1 _6048_ (.A(_1694_),
    .B(net359),
    .Y(_3060_));
 sky130_fd_sc_hd__nand2_1 _6049_ (.A(_1697_),
    .B(_3060_),
    .Y(_3061_));
 sky130_fd_sc_hd__nor2_1 _6050_ (.A(_1697_),
    .B(_3060_),
    .Y(_3062_));
 sky130_fd_sc_hd__or2_1 _6051_ (.A(_1697_),
    .B(_3060_),
    .X(_3063_));
 sky130_fd_sc_hd__nand2_1 _6052_ (.A(_3061_),
    .B(_3063_),
    .Y(_3064_));
 sky130_fd_sc_hd__o21ai_1 _6053_ (.A1(_3059_),
    .A2(_3064_),
    .B1(net317),
    .Y(_3065_));
 sky130_fd_sc_hd__a21o_1 _6054_ (.A1(_3059_),
    .A2(_3064_),
    .B1(_3065_),
    .X(_3066_));
 sky130_fd_sc_hd__mux4_1 _6055_ (.A0(_1638_),
    .A1(_1697_),
    .A2(_1629_),
    .A3(_1660_),
    .S0(net200),
    .S1(net194),
    .X(_3067_));
 sky130_fd_sc_hd__mux2_1 _6056_ (.A0(_2983_),
    .A1(_3067_),
    .S(net206),
    .X(_3068_));
 sky130_fd_sc_hd__or2_1 _6057_ (.A(net209),
    .B(_3068_),
    .X(_3069_));
 sky130_fd_sc_hd__o21ai_1 _6058_ (.A1(net213),
    .A2(_2883_),
    .B1(_3069_),
    .Y(_3070_));
 sky130_fd_sc_hd__mux2_1 _6059_ (.A0(_2872_),
    .A1(_2877_),
    .S(net213),
    .X(_3071_));
 sky130_fd_sc_hd__a2bb2o_2 _6060_ (.A1_N(_2721_),
    .A2_N(_3070_),
    .B1(_3071_),
    .B2(_2691_),
    .X(_3072_));
 sky130_fd_sc_hd__a221o_1 _6061_ (.A1(_1694_),
    .A2(net360),
    .B1(net357),
    .B2(_1698_),
    .C1(net362),
    .X(_3073_));
 sky130_fd_sc_hd__o21a_1 _6062_ (.A1(_2835_),
    .A2(_2873_),
    .B1(net211),
    .X(_3074_));
 sky130_fd_sc_hd__nor2_1 _6063_ (.A(_2989_),
    .B(_3074_),
    .Y(_3075_));
 sky130_fd_sc_hd__a2bb2o_2 _6064_ (.A1_N(_2687_),
    .A2_N(_3075_),
    .B1(_2940_),
    .B2(_2873_),
    .X(_3076_));
 sky130_fd_sc_hd__a221o_1 _6065_ (.A1(_1699_),
    .A2(_3073_),
    .B1(_3076_),
    .B2(net187),
    .C1(net223),
    .X(_3077_));
 sky130_fd_sc_hd__a21oi_1 _6066_ (.A1(net190),
    .A2(_3072_),
    .B1(_3077_),
    .Y(_3078_));
 sky130_fd_sc_hd__a221oi_1 _6067_ (.A1(net2289),
    .A2(net223),
    .B1(_3066_),
    .B2(_3078_),
    .C1(net467),
    .Y(_0729_));
 sky130_fd_sc_hd__xnor2_1 _6068_ (.A(_1670_),
    .B(net359),
    .Y(_3079_));
 sky130_fd_sc_hd__and2_1 _6069_ (.A(_1673_),
    .B(_3079_),
    .X(_3080_));
 sky130_fd_sc_hd__nand2_1 _6070_ (.A(_1673_),
    .B(_3079_),
    .Y(_3081_));
 sky130_fd_sc_hd__nor2_1 _6071_ (.A(_1673_),
    .B(_3079_),
    .Y(_3082_));
 sky130_fd_sc_hd__nor2_1 _6072_ (.A(_3080_),
    .B(_3082_),
    .Y(_3083_));
 sky130_fd_sc_hd__a21o_1 _6073_ (.A1(_3059_),
    .A2(_3061_),
    .B1(_3062_),
    .X(_3084_));
 sky130_fd_sc_hd__nand2_1 _6074_ (.A(_3083_),
    .B(_3084_),
    .Y(_3085_));
 sky130_fd_sc_hd__or2_1 _6075_ (.A(_3083_),
    .B(_3084_),
    .X(_3086_));
 sky130_fd_sc_hd__a21oi_1 _6076_ (.A1(_3085_),
    .A2(_3086_),
    .B1(_2731_),
    .Y(_3087_));
 sky130_fd_sc_hd__mux4_1 _6077_ (.A0(_1660_),
    .A1(_1673_),
    .A2(_1638_),
    .A3(_1697_),
    .S0(net200),
    .S1(net192),
    .X(_3088_));
 sky130_fd_sc_hd__inv_2 _6078_ (.A(_3088_),
    .Y(_3089_));
 sky130_fd_sc_hd__mux2_1 _6079_ (.A0(_3007_),
    .A1(_3089_),
    .S(net206),
    .X(_3090_));
 sky130_fd_sc_hd__mux2_1 _6080_ (.A0(_2910_),
    .A1(_3090_),
    .S(net213),
    .X(_3091_));
 sky130_fd_sc_hd__or2_1 _6081_ (.A(_2721_),
    .B(_3091_),
    .X(_3092_));
 sky130_fd_sc_hd__mux2_1 _6082_ (.A0(_2896_),
    .A1(_2912_),
    .S(net213),
    .X(_3093_));
 sky130_fd_sc_hd__a21bo_1 _6083_ (.A1(_2691_),
    .A2(_3093_),
    .B1_N(_3092_),
    .X(_3094_));
 sky130_fd_sc_hd__a221o_1 _6084_ (.A1(_1674_),
    .A2(net362),
    .B1(net360),
    .B2(_1670_),
    .C1(net224),
    .X(_3095_));
 sky130_fd_sc_hd__a22o_1 _6085_ (.A1(net357),
    .A2(_3083_),
    .B1(_3094_),
    .B2(net190),
    .X(_3096_));
 sky130_fd_sc_hd__o21ba_1 _6086_ (.A1(net207),
    .A2(_2901_),
    .B1_N(_2989_),
    .X(_3097_));
 sky130_fd_sc_hd__a2bb2o_2 _6087_ (.A1_N(_2687_),
    .A2_N(_3097_),
    .B1(_2940_),
    .B2(_2898_),
    .X(_3098_));
 sky130_fd_sc_hd__a211o_1 _6088_ (.A1(net186),
    .A2(_3098_),
    .B1(_3096_),
    .C1(_3095_),
    .X(_3099_));
 sky130_fd_sc_hd__a21o_1 _6089_ (.A1(_1670_),
    .A2(_1673_),
    .B1(_2737_),
    .X(_3100_));
 sky130_fd_sc_hd__o211a_1 _6090_ (.A1(_3087_),
    .A2(_3099_),
    .B1(_3100_),
    .C1(net443),
    .X(_0730_));
 sky130_fd_sc_hd__a21o_1 _6091_ (.A1(_3081_),
    .A2(_3084_),
    .B1(_3082_),
    .X(_3101_));
 sky130_fd_sc_hd__xnor2_1 _6092_ (.A(_1682_),
    .B(net359),
    .Y(_3102_));
 sky130_fd_sc_hd__nand2_1 _6093_ (.A(_1684_),
    .B(_3102_),
    .Y(_3103_));
 sky130_fd_sc_hd__or2_1 _6094_ (.A(_1684_),
    .B(_3102_),
    .X(_3104_));
 sky130_fd_sc_hd__nand2_1 _6095_ (.A(_3103_),
    .B(_3104_),
    .Y(_3105_));
 sky130_fd_sc_hd__nor2_1 _6096_ (.A(_3101_),
    .B(_3105_),
    .Y(_3106_));
 sky130_fd_sc_hd__a21o_1 _6097_ (.A1(_3101_),
    .A2(_3105_),
    .B1(_2731_),
    .X(_3107_));
 sky130_fd_sc_hd__mux4_1 _6098_ (.A0(_1684_),
    .A1(_1697_),
    .A2(_1673_),
    .A3(_1660_),
    .S0(net197),
    .S1(net192),
    .X(_3108_));
 sky130_fd_sc_hd__mux2_1 _6099_ (.A0(_3026_),
    .A1(_3108_),
    .S(net205),
    .X(_3109_));
 sky130_fd_sc_hd__nor2_1 _6100_ (.A(net207),
    .B(_3109_),
    .Y(_3110_));
 sky130_fd_sc_hd__a211o_1 _6101_ (.A1(net207),
    .A2(_2934_),
    .B1(_3110_),
    .C1(_2721_),
    .X(_3111_));
 sky130_fd_sc_hd__mux2_1 _6102_ (.A0(_2929_),
    .A1(_2936_),
    .S(net207),
    .X(_3112_));
 sky130_fd_sc_hd__a21boi_2 _6103_ (.A1(_2691_),
    .A2(_3112_),
    .B1_N(_3111_),
    .Y(_3113_));
 sky130_fd_sc_hd__a221o_1 _6104_ (.A1(_1682_),
    .A2(net360),
    .B1(net357),
    .B2(_1685_),
    .C1(net362),
    .X(_3114_));
 sky130_fd_sc_hd__o21ai_1 _6105_ (.A1(_1682_),
    .A2(_1684_),
    .B1(_3114_),
    .Y(_3115_));
 sky130_fd_sc_hd__a21oi_1 _6106_ (.A1(net211),
    .A2(_2938_),
    .B1(_2989_),
    .Y(_3116_));
 sky130_fd_sc_hd__o32a_4 _6107_ (.A1(net207),
    .A2(_2689_),
    .A3(_2943_),
    .B1(_3116_),
    .B2(_2687_),
    .X(_3117_));
 sky130_fd_sc_hd__o211a_1 _6108_ (.A1(net187),
    .A2(_3113_),
    .B1(_3115_),
    .C1(_2737_),
    .X(_3118_));
 sky130_fd_sc_hd__o22a_1 _6109_ (.A1(_3106_),
    .A2(_3107_),
    .B1(_3117_),
    .B2(net190),
    .X(_3119_));
 sky130_fd_sc_hd__a221oi_2 _6110_ (.A1(_1685_),
    .A2(net224),
    .B1(_3118_),
    .B2(_3119_),
    .C1(net467),
    .Y(_0731_));
 sky130_fd_sc_hd__xnor2_1 _6111_ (.A(_1705_),
    .B(net359),
    .Y(_3120_));
 sky130_fd_sc_hd__and2_1 _6112_ (.A(_1707_),
    .B(_3120_),
    .X(_3121_));
 sky130_fd_sc_hd__nand2_1 _6113_ (.A(_1707_),
    .B(_3120_),
    .Y(_3122_));
 sky130_fd_sc_hd__nor2_1 _6114_ (.A(_1707_),
    .B(_3120_),
    .Y(_3123_));
 sky130_fd_sc_hd__nor2_1 _6115_ (.A(_3121_),
    .B(_3123_),
    .Y(_3124_));
 sky130_fd_sc_hd__a21bo_1 _6116_ (.A1(_3101_),
    .A2(_3103_),
    .B1_N(_3104_),
    .X(_3125_));
 sky130_fd_sc_hd__xnor2_1 _6117_ (.A(_3124_),
    .B(_3125_),
    .Y(_3126_));
 sky130_fd_sc_hd__mux4_1 _6118_ (.A0(_1673_),
    .A1(_1697_),
    .A2(_1707_),
    .A3(_1684_),
    .S0(net192),
    .S1(net199),
    .X(_3127_));
 sky130_fd_sc_hd__mux2_1 _6119_ (.A0(_3046_),
    .A1(_3127_),
    .S(net205),
    .X(_3128_));
 sky130_fd_sc_hd__mux2_4 _6120_ (.A0(_2958_),
    .A1(_3128_),
    .S(net212),
    .X(_3129_));
 sky130_fd_sc_hd__a221o_1 _6121_ (.A1(_1708_),
    .A2(net362),
    .B1(net360),
    .B2(_1705_),
    .C1(net223),
    .X(_3130_));
 sky130_fd_sc_hd__a221o_1 _6122_ (.A1(net357),
    .A2(_3124_),
    .B1(_3129_),
    .B2(_2722_),
    .C1(_3130_),
    .X(_3131_));
 sky130_fd_sc_hd__o21a_4 _6123_ (.A1(_1337_),
    .A2(net188),
    .B1(_2686_),
    .X(_3132_));
 sky130_fd_sc_hd__o21ai_4 _6124_ (.A1(_1337_),
    .A2(net188),
    .B1(_2686_),
    .Y(_3133_));
 sky130_fd_sc_hd__nand2_1 _6125_ (.A(net212),
    .B(_2970_),
    .Y(_3134_));
 sky130_fd_sc_hd__a21oi_1 _6126_ (.A1(net185),
    .A2(_3134_),
    .B1(_2689_),
    .Y(_3135_));
 sky130_fd_sc_hd__mux2_1 _6127_ (.A0(_2961_),
    .A1(_2968_),
    .S(net207),
    .X(_3136_));
 sky130_fd_sc_hd__o22a_1 _6128_ (.A1(_3132_),
    .A2(_3135_),
    .B1(_3136_),
    .B2(net184),
    .X(_3137_));
 sky130_fd_sc_hd__a211o_1 _6129_ (.A1(net317),
    .A2(_3126_),
    .B1(_3131_),
    .C1(_3137_),
    .X(_3138_));
 sky130_fd_sc_hd__a21o_1 _6130_ (.A1(_1705_),
    .A2(_1707_),
    .B1(_2737_),
    .X(_3139_));
 sky130_fd_sc_hd__and3_2 _6131_ (.A(net443),
    .B(_3138_),
    .C(_3139_),
    .X(_0732_));
 sky130_fd_sc_hd__a21o_1 _6132_ (.A1(_3122_),
    .A2(_3125_),
    .B1(_3123_),
    .X(_3140_));
 sky130_fd_sc_hd__xnor2_1 _6133_ (.A(_1411_),
    .B(_2729_),
    .Y(_3141_));
 sky130_fd_sc_hd__nand2_1 _6134_ (.A(_1414_),
    .B(_3141_),
    .Y(_3142_));
 sky130_fd_sc_hd__nor2_1 _6135_ (.A(_1414_),
    .B(_3141_),
    .Y(_3143_));
 sky130_fd_sc_hd__inv_2 _6136_ (.A(_3143_),
    .Y(_3144_));
 sky130_fd_sc_hd__a21bo_1 _6137_ (.A1(_3142_),
    .A2(_3144_),
    .B1_N(_3140_),
    .X(_3145_));
 sky130_fd_sc_hd__or3b_1 _6138_ (.A(_3143_),
    .B(_3140_),
    .C_N(_3142_),
    .X(_3146_));
 sky130_fd_sc_hd__mux4_1 _6139_ (.A0(_1414_),
    .A1(_1684_),
    .A2(_1707_),
    .A3(_1673_),
    .S0(net198),
    .S1(net194),
    .X(_3147_));
 sky130_fd_sc_hd__mux2_1 _6140_ (.A0(_3067_),
    .A1(_3147_),
    .S(net206),
    .X(_3148_));
 sky130_fd_sc_hd__mux2_1 _6141_ (.A0(_2984_),
    .A1(_3148_),
    .S(net213),
    .X(_3149_));
 sky130_fd_sc_hd__nand2_1 _6142_ (.A(net186),
    .B(_2719_),
    .Y(_3150_));
 sky130_fd_sc_hd__o211a_1 _6143_ (.A1(net186),
    .A2(_3149_),
    .B1(_3150_),
    .C1(_2720_),
    .X(_3151_));
 sky130_fd_sc_hd__nor2_4 _6144_ (.A(net184),
    .B(_2689_),
    .Y(_3152_));
 sky130_fd_sc_hd__a221o_1 _6145_ (.A1(_1412_),
    .A2(net360),
    .B1(net357),
    .B2(_1415_),
    .C1(net362),
    .X(_3153_));
 sky130_fd_sc_hd__o21a_1 _6146_ (.A1(_1412_),
    .A2(_1414_),
    .B1(_3153_),
    .X(_3154_));
 sky130_fd_sc_hd__o21a_1 _6147_ (.A1(net186),
    .A2(_2716_),
    .B1(_3132_),
    .X(_3155_));
 sky130_fd_sc_hd__a2111o_1 _6148_ (.A1(_2716_),
    .A2(_3152_),
    .B1(_3154_),
    .C1(_3155_),
    .D1(net223),
    .X(_3156_));
 sky130_fd_sc_hd__a311o_1 _6149_ (.A1(net317),
    .A2(_3145_),
    .A3(_3146_),
    .B1(_3151_),
    .C1(_3156_),
    .X(_3157_));
 sky130_fd_sc_hd__nand2_1 _6150_ (.A(_1415_),
    .B(net224),
    .Y(_3158_));
 sky130_fd_sc_hd__and3_1 _6151_ (.A(net444),
    .B(_3157_),
    .C(_3158_),
    .X(_0733_));
 sky130_fd_sc_hd__xnor2_1 _6152_ (.A(_1388_),
    .B(net359),
    .Y(_3159_));
 sky130_fd_sc_hd__nand2_1 _6153_ (.A(_1391_),
    .B(_3159_),
    .Y(_3160_));
 sky130_fd_sc_hd__nor2_1 _6154_ (.A(_1391_),
    .B(_3159_),
    .Y(_3161_));
 sky130_fd_sc_hd__xnor2_1 _6155_ (.A(_1390_),
    .B(_3159_),
    .Y(_3162_));
 sky130_fd_sc_hd__a21o_1 _6156_ (.A1(_3140_),
    .A2(_3142_),
    .B1(_3143_),
    .X(_3163_));
 sky130_fd_sc_hd__xnor2_1 _6157_ (.A(_3162_),
    .B(_3163_),
    .Y(_3164_));
 sky130_fd_sc_hd__mux4_1 _6158_ (.A0(_1391_),
    .A1(_1414_),
    .A2(_1707_),
    .A3(_1684_),
    .S0(net193),
    .S1(net197),
    .X(_3165_));
 sky130_fd_sc_hd__mux2_1 _6159_ (.A0(_3088_),
    .A1(_3165_),
    .S(net206),
    .X(_3166_));
 sky130_fd_sc_hd__mux2_1 _6160_ (.A0(_3008_),
    .A1(_3166_),
    .S(net214),
    .X(_3167_));
 sky130_fd_sc_hd__nand2_1 _6161_ (.A(net186),
    .B(_2776_),
    .Y(_3168_));
 sky130_fd_sc_hd__o211a_1 _6162_ (.A1(net186),
    .A2(_3167_),
    .B1(_3168_),
    .C1(_2720_),
    .X(_3169_));
 sky130_fd_sc_hd__a221o_1 _6163_ (.A1(_1392_),
    .A2(net362),
    .B1(_2727_),
    .B2(_1388_),
    .C1(net224),
    .X(_3170_));
 sky130_fd_sc_hd__a221o_1 _6164_ (.A1(_2762_),
    .A2(_3152_),
    .B1(_3162_),
    .B2(net357),
    .C1(_3170_),
    .X(_3171_));
 sky130_fd_sc_hd__or2_1 _6165_ (.A(net186),
    .B(_2758_),
    .X(_3172_));
 sky130_fd_sc_hd__a221o_1 _6166_ (.A1(net317),
    .A2(_3164_),
    .B1(_3172_),
    .B2(_3132_),
    .C1(_3171_),
    .X(_3173_));
 sky130_fd_sc_hd__nand2_1 _6167_ (.A(_1393_),
    .B(net223),
    .Y(_3174_));
 sky130_fd_sc_hd__o211a_1 _6168_ (.A1(_3169_),
    .A2(_3173_),
    .B1(_3174_),
    .C1(net444),
    .X(_0734_));
 sky130_fd_sc_hd__a21o_1 _6169_ (.A1(_3160_),
    .A2(_3163_),
    .B1(_3161_),
    .X(_3175_));
 sky130_fd_sc_hd__xnor2_1 _6170_ (.A(_1423_),
    .B(net359),
    .Y(_3176_));
 sky130_fd_sc_hd__nand2_1 _6171_ (.A(_1425_),
    .B(_3176_),
    .Y(_3177_));
 sky130_fd_sc_hd__nor2_1 _6172_ (.A(_1425_),
    .B(_3176_),
    .Y(_3178_));
 sky130_fd_sc_hd__inv_2 _6173_ (.A(_3178_),
    .Y(_3179_));
 sky130_fd_sc_hd__or3b_1 _6174_ (.A(_3178_),
    .B(_3175_),
    .C_N(_3177_),
    .X(_3180_));
 sky130_fd_sc_hd__a21bo_1 _6175_ (.A1(_3177_),
    .A2(_3179_),
    .B1_N(_3175_),
    .X(_3181_));
 sky130_fd_sc_hd__a2111oi_2 _6176_ (.A1(_1338_),
    .A2(net184),
    .B1(_2687_),
    .C1(_2812_),
    .D1(_2816_),
    .Y(_3182_));
 sky130_fd_sc_hd__a221o_1 _6177_ (.A1(_1423_),
    .A2(net360),
    .B1(net357),
    .B2(_1426_),
    .C1(net362),
    .X(_3183_));
 sky130_fd_sc_hd__a32o_2 _6178_ (.A1(net212),
    .A2(_2720_),
    .A3(_2794_),
    .B1(_2686_),
    .B2(_1337_),
    .X(_3184_));
 sky130_fd_sc_hd__a221o_1 _6179_ (.A1(_1427_),
    .A2(_3183_),
    .B1(_3184_),
    .B2(net186),
    .C1(net223),
    .X(_3185_));
 sky130_fd_sc_hd__mux4_1 _6180_ (.A0(_1414_),
    .A1(_1707_),
    .A2(_1425_),
    .A3(_1391_),
    .S0(net193),
    .S1(net199),
    .X(_3186_));
 sky130_fd_sc_hd__mux2_1 _6181_ (.A0(_3108_),
    .A1(_3186_),
    .S(net205),
    .X(_3187_));
 sky130_fd_sc_hd__mux2_1 _6182_ (.A0(_3027_),
    .A1(_3187_),
    .S(net212),
    .X(_3188_));
 sky130_fd_sc_hd__a21bo_1 _6183_ (.A1(_2720_),
    .A2(_3188_),
    .B1_N(_2813_),
    .X(_3189_));
 sky130_fd_sc_hd__a32o_1 _6184_ (.A1(_2732_),
    .A2(_3180_),
    .A3(_3181_),
    .B1(_3189_),
    .B2(net190),
    .X(_3190_));
 sky130_fd_sc_hd__a21oi_1 _6185_ (.A1(_1426_),
    .A2(net223),
    .B1(net467),
    .Y(_3191_));
 sky130_fd_sc_hd__o31a_2 _6186_ (.A1(_3182_),
    .A2(_3185_),
    .A3(_3190_),
    .B1(_3191_),
    .X(_0735_));
 sky130_fd_sc_hd__xnor2_1 _6187_ (.A(_1399_),
    .B(net359),
    .Y(_3192_));
 sky130_fd_sc_hd__and2_1 _6188_ (.A(_1401_),
    .B(_3192_),
    .X(_3193_));
 sky130_fd_sc_hd__nand2_1 _6189_ (.A(_1401_),
    .B(_3192_),
    .Y(_3194_));
 sky130_fd_sc_hd__nor2_1 _6190_ (.A(_1401_),
    .B(_3192_),
    .Y(_3195_));
 sky130_fd_sc_hd__nor2_1 _6191_ (.A(_3193_),
    .B(_3195_),
    .Y(_3196_));
 sky130_fd_sc_hd__a21o_1 _6192_ (.A1(_3175_),
    .A2(_3177_),
    .B1(_3178_),
    .X(_3197_));
 sky130_fd_sc_hd__xnor2_1 _6193_ (.A(_3196_),
    .B(_3197_),
    .Y(_3198_));
 sky130_fd_sc_hd__mux4_1 _6194_ (.A0(_1391_),
    .A1(_1401_),
    .A2(_1414_),
    .A3(_1425_),
    .S0(net199),
    .S1(net193),
    .X(_3199_));
 sky130_fd_sc_hd__mux2_1 _6195_ (.A0(_3127_),
    .A1(_3199_),
    .S(net205),
    .X(_3200_));
 sky130_fd_sc_hd__mux2_1 _6196_ (.A0(_3047_),
    .A1(_3200_),
    .S(net214),
    .X(_3201_));
 sky130_fd_sc_hd__or2_1 _6197_ (.A(net190),
    .B(_2851_),
    .X(_3202_));
 sky130_fd_sc_hd__o211a_1 _6198_ (.A1(net186),
    .A2(_3201_),
    .B1(_3202_),
    .C1(_2720_),
    .X(_3203_));
 sky130_fd_sc_hd__a221o_1 _6199_ (.A1(_1402_),
    .A2(net362),
    .B1(net360),
    .B2(_1399_),
    .C1(net223),
    .X(_3204_));
 sky130_fd_sc_hd__a221o_1 _6200_ (.A1(_2840_),
    .A2(_3152_),
    .B1(_3196_),
    .B2(net357),
    .C1(_3204_),
    .X(_3205_));
 sky130_fd_sc_hd__or2_1 _6201_ (.A(net186),
    .B(_2837_),
    .X(_3206_));
 sky130_fd_sc_hd__a221o_1 _6202_ (.A1(_2732_),
    .A2(_3198_),
    .B1(_3206_),
    .B2(_3132_),
    .C1(_3205_),
    .X(_3207_));
 sky130_fd_sc_hd__a21o_1 _6203_ (.A1(_1399_),
    .A2(_1401_),
    .B1(_2737_),
    .X(_3208_));
 sky130_fd_sc_hd__o211a_1 _6204_ (.A1(_3203_),
    .A2(_3207_),
    .B1(_3208_),
    .C1(net444),
    .X(_0736_));
 sky130_fd_sc_hd__a21o_1 _6205_ (.A1(_3194_),
    .A2(_3197_),
    .B1(_3195_),
    .X(_3209_));
 sky130_fd_sc_hd__xnor2_1 _6206_ (.A(_1456_),
    .B(net359),
    .Y(_3210_));
 sky130_fd_sc_hd__nand2_1 _6207_ (.A(_1458_),
    .B(_3210_),
    .Y(_3211_));
 sky130_fd_sc_hd__nor2_1 _6208_ (.A(_1458_),
    .B(_3210_),
    .Y(_3212_));
 sky130_fd_sc_hd__or2_1 _6209_ (.A(_1458_),
    .B(_3210_),
    .X(_3213_));
 sky130_fd_sc_hd__nand2_1 _6210_ (.A(_3211_),
    .B(_3213_),
    .Y(_3214_));
 sky130_fd_sc_hd__nand2_1 _6211_ (.A(_3209_),
    .B(_3214_),
    .Y(_3215_));
 sky130_fd_sc_hd__or2_1 _6212_ (.A(_3209_),
    .B(_3214_),
    .X(_3216_));
 sky130_fd_sc_hd__mux4_1 _6213_ (.A0(_1458_),
    .A1(_1425_),
    .A2(_1401_),
    .A3(_1391_),
    .S0(net198),
    .S1(net194),
    .X(_3217_));
 sky130_fd_sc_hd__mux2_1 _6214_ (.A0(_3147_),
    .A1(_3217_),
    .S(net206),
    .X(_3218_));
 sky130_fd_sc_hd__o31a_1 _6215_ (.A1(net209),
    .A2(net186),
    .A3(_3218_),
    .B1(_2720_),
    .X(_3219_));
 sky130_fd_sc_hd__o221a_1 _6216_ (.A1(net190),
    .A2(_2885_),
    .B1(_3068_),
    .B2(net213),
    .C1(_3219_),
    .X(_3220_));
 sky130_fd_sc_hd__o21a_1 _6217_ (.A1(net211),
    .A2(_2873_),
    .B1(_3152_),
    .X(_3221_));
 sky130_fd_sc_hd__o22a_1 _6218_ (.A1(net184),
    .A2(_2875_),
    .B1(_3132_),
    .B2(_3221_),
    .X(_3222_));
 sky130_fd_sc_hd__a221o_1 _6219_ (.A1(_1456_),
    .A2(net360),
    .B1(net356),
    .B2(_1459_),
    .C1(net362),
    .X(_3223_));
 sky130_fd_sc_hd__o21a_1 _6220_ (.A1(_1456_),
    .A2(_1458_),
    .B1(_3223_),
    .X(_3224_));
 sky130_fd_sc_hd__or4_1 _6221_ (.A(net223),
    .B(_3220_),
    .C(_3222_),
    .D(_3224_),
    .X(_3225_));
 sky130_fd_sc_hd__a31o_1 _6222_ (.A1(net317),
    .A2(_3215_),
    .A3(_3216_),
    .B1(_3225_),
    .X(_3226_));
 sky130_fd_sc_hd__nand2_1 _6223_ (.A(_1459_),
    .B(net223),
    .Y(_3227_));
 sky130_fd_sc_hd__and3_1 _6224_ (.A(net438),
    .B(_3226_),
    .C(_3227_),
    .X(_0737_));
 sky130_fd_sc_hd__xnor2_1 _6225_ (.A(_1435_),
    .B(net358),
    .Y(_3228_));
 sky130_fd_sc_hd__and2_1 _6226_ (.A(_1437_),
    .B(_3228_),
    .X(_3229_));
 sky130_fd_sc_hd__nand2_1 _6227_ (.A(_1437_),
    .B(_3228_),
    .Y(_3230_));
 sky130_fd_sc_hd__nor2_1 _6228_ (.A(_1437_),
    .B(_3228_),
    .Y(_3231_));
 sky130_fd_sc_hd__nor2_1 _6229_ (.A(_3229_),
    .B(_3231_),
    .Y(_3232_));
 sky130_fd_sc_hd__a21o_1 _6230_ (.A1(_3209_),
    .A2(_3211_),
    .B1(_3212_),
    .X(_3233_));
 sky130_fd_sc_hd__xor2_1 _6231_ (.A(_3232_),
    .B(_3233_),
    .X(_3234_));
 sky130_fd_sc_hd__o21ai_1 _6232_ (.A1(net185),
    .A2(_2902_),
    .B1(_3132_),
    .Y(_3235_));
 sky130_fd_sc_hd__a221o_1 _6233_ (.A1(_1438_),
    .A2(net363),
    .B1(net361),
    .B2(_1435_),
    .C1(net222),
    .X(_3236_));
 sky130_fd_sc_hd__a21oi_1 _6234_ (.A1(net356),
    .A2(_3232_),
    .B1(_3236_),
    .Y(_3237_));
 sky130_fd_sc_hd__mux4_1 _6235_ (.A0(_1401_),
    .A1(_1425_),
    .A2(_1437_),
    .A3(_1458_),
    .S0(net193),
    .S1(net200),
    .X(_3238_));
 sky130_fd_sc_hd__mux2_1 _6236_ (.A0(_3165_),
    .A1(_3238_),
    .S(net206),
    .X(_3239_));
 sky130_fd_sc_hd__nand2_1 _6237_ (.A(net213),
    .B(_3239_),
    .Y(_3240_));
 sky130_fd_sc_hd__o211a_1 _6238_ (.A1(net213),
    .A2(_3090_),
    .B1(_3240_),
    .C1(net188),
    .X(_3241_));
 sky130_fd_sc_hd__o31a_1 _6239_ (.A1(net209),
    .A2(_2721_),
    .A3(_2910_),
    .B1(_2723_),
    .X(_3242_));
 sky130_fd_sc_hd__o22a_1 _6240_ (.A1(_2731_),
    .A2(_3234_),
    .B1(_3241_),
    .B2(_3242_),
    .X(_3243_));
 sky130_fd_sc_hd__o211a_1 _6241_ (.A1(net185),
    .A2(_2900_),
    .B1(_3237_),
    .C1(_3243_),
    .X(_3244_));
 sky130_fd_sc_hd__a21oi_1 _6242_ (.A1(_1435_),
    .A2(_1437_),
    .B1(net221),
    .Y(_3245_));
 sky130_fd_sc_hd__a211oi_1 _6243_ (.A1(_3235_),
    .A2(_3244_),
    .B1(_3245_),
    .C1(net467),
    .Y(_0738_));
 sky130_fd_sc_hd__a21o_1 _6244_ (.A1(_3230_),
    .A2(_3233_),
    .B1(_3231_),
    .X(_3246_));
 sky130_fd_sc_hd__xnor2_1 _6245_ (.A(_1445_),
    .B(net358),
    .Y(_3247_));
 sky130_fd_sc_hd__nand2_1 _6246_ (.A(_1447_),
    .B(_3247_),
    .Y(_3248_));
 sky130_fd_sc_hd__nor2_1 _6247_ (.A(_1447_),
    .B(_3247_),
    .Y(_3249_));
 sky130_fd_sc_hd__inv_2 _6248_ (.A(_3249_),
    .Y(_3250_));
 sky130_fd_sc_hd__a21oi_1 _6249_ (.A1(_3248_),
    .A2(_3250_),
    .B1(_3246_),
    .Y(_3251_));
 sky130_fd_sc_hd__and3_1 _6250_ (.A(_3246_),
    .B(_3248_),
    .C(_3250_),
    .X(_3252_));
 sky130_fd_sc_hd__o21a_1 _6251_ (.A1(_3251_),
    .A2(_3252_),
    .B1(net317),
    .X(_3253_));
 sky130_fd_sc_hd__mux4_1 _6252_ (.A0(_1447_),
    .A1(_1458_),
    .A2(_1437_),
    .A3(_1401_),
    .S0(net197),
    .S1(net193),
    .X(_3254_));
 sky130_fd_sc_hd__mux2_1 _6253_ (.A0(_3186_),
    .A1(_3254_),
    .S(net204),
    .X(_3255_));
 sky130_fd_sc_hd__mux2_1 _6254_ (.A0(_3109_),
    .A1(_3255_),
    .S(net212),
    .X(_3256_));
 sky130_fd_sc_hd__o2bb2a_1 _6255_ (.A1_N(_2723_),
    .A2_N(_2935_),
    .B1(_3256_),
    .B2(net184),
    .X(_3257_));
 sky130_fd_sc_hd__a221o_1 _6256_ (.A1(_1445_),
    .A2(net361),
    .B1(net356),
    .B2(_1448_),
    .C1(net363),
    .X(_3258_));
 sky130_fd_sc_hd__o21a_1 _6257_ (.A1(_1445_),
    .A2(_1447_),
    .B1(_3258_),
    .X(_3259_));
 sky130_fd_sc_hd__a21oi_1 _6258_ (.A1(net188),
    .A2(_2939_),
    .B1(_3133_),
    .Y(_3260_));
 sky130_fd_sc_hd__a2111o_1 _6259_ (.A1(net188),
    .A2(_2944_),
    .B1(_3257_),
    .C1(_3259_),
    .D1(net224),
    .X(_3261_));
 sky130_fd_sc_hd__nand2_1 _6260_ (.A(net2295),
    .B(net224),
    .Y(_3262_));
 sky130_fd_sc_hd__o311a_1 _6261_ (.A1(_3253_),
    .A2(_3260_),
    .A3(_3261_),
    .B1(_3262_),
    .C1(net438),
    .X(_0739_));
 sky130_fd_sc_hd__xnor2_1 _6262_ (.A(_1466_),
    .B(net358),
    .Y(_3263_));
 sky130_fd_sc_hd__and2_1 _6263_ (.A(_1468_),
    .B(_3263_),
    .X(_3264_));
 sky130_fd_sc_hd__nand2_1 _6264_ (.A(_1468_),
    .B(_3263_),
    .Y(_3265_));
 sky130_fd_sc_hd__nor2_1 _6265_ (.A(_1468_),
    .B(_3263_),
    .Y(_3266_));
 sky130_fd_sc_hd__nor2_1 _6266_ (.A(_3264_),
    .B(_3266_),
    .Y(_3267_));
 sky130_fd_sc_hd__a21o_1 _6267_ (.A1(_3246_),
    .A2(_3248_),
    .B1(_3249_),
    .X(_3268_));
 sky130_fd_sc_hd__xnor2_1 _6268_ (.A(_3267_),
    .B(_3268_),
    .Y(_3269_));
 sky130_fd_sc_hd__a21oi_1 _6269_ (.A1(net188),
    .A2(_2972_),
    .B1(_3133_),
    .Y(_3270_));
 sky130_fd_sc_hd__a221o_1 _6270_ (.A1(_1469_),
    .A2(net363),
    .B1(net361),
    .B2(_1466_),
    .C1(net222),
    .X(_3271_));
 sky130_fd_sc_hd__a221o_1 _6271_ (.A1(net188),
    .A2(_2971_),
    .B1(_3267_),
    .B2(net356),
    .C1(_3271_),
    .X(_3272_));
 sky130_fd_sc_hd__mux4_1 _6272_ (.A0(_1437_),
    .A1(_1458_),
    .A2(_1468_),
    .A3(_1447_),
    .S0(net193),
    .S1(net199),
    .X(_3273_));
 sky130_fd_sc_hd__mux2_1 _6273_ (.A0(_3199_),
    .A1(_3273_),
    .S(net204),
    .X(_3274_));
 sky130_fd_sc_hd__mux2_1 _6274_ (.A0(_3128_),
    .A1(_3274_),
    .S(net212),
    .X(_3275_));
 sky130_fd_sc_hd__o22a_1 _6275_ (.A1(_2722_),
    .A2(_2959_),
    .B1(_3275_),
    .B2(net185),
    .X(_3276_));
 sky130_fd_sc_hd__a211o_1 _6276_ (.A1(net317),
    .A2(_3269_),
    .B1(_3272_),
    .C1(_3276_),
    .X(_3277_));
 sky130_fd_sc_hd__a21o_1 _6277_ (.A1(_1466_),
    .A2(_1468_),
    .B1(net221),
    .X(_3278_));
 sky130_fd_sc_hd__o211a_1 _6278_ (.A1(_3270_),
    .A2(_3277_),
    .B1(_3278_),
    .C1(net438),
    .X(_0740_));
 sky130_fd_sc_hd__a21o_1 _6279_ (.A1(_3265_),
    .A2(_3268_),
    .B1(_3266_),
    .X(_3279_));
 sky130_fd_sc_hd__xnor2_1 _6280_ (.A(_1502_),
    .B(net358),
    .Y(_3280_));
 sky130_fd_sc_hd__nand2_1 _6281_ (.A(_1505_),
    .B(_3280_),
    .Y(_3281_));
 sky130_fd_sc_hd__nor2_1 _6282_ (.A(_1505_),
    .B(_3280_),
    .Y(_3282_));
 sky130_fd_sc_hd__inv_2 _6283_ (.A(_3282_),
    .Y(_3283_));
 sky130_fd_sc_hd__a21oi_1 _6284_ (.A1(_3281_),
    .A2(_3283_),
    .B1(_3279_),
    .Y(_3284_));
 sky130_fd_sc_hd__and3_1 _6285_ (.A(_3279_),
    .B(_3281_),
    .C(_3283_),
    .X(_3285_));
 sky130_fd_sc_hd__o21a_1 _6286_ (.A1(_3284_),
    .A2(_3285_),
    .B1(net317),
    .X(_3286_));
 sky130_fd_sc_hd__mux4_1 _6287_ (.A0(_1447_),
    .A1(_1505_),
    .A2(_1437_),
    .A3(_1468_),
    .S0(net199),
    .S1(net193),
    .X(_3287_));
 sky130_fd_sc_hd__mux2_1 _6288_ (.A0(_3217_),
    .A1(_3287_),
    .S(net206),
    .X(_3288_));
 sky130_fd_sc_hd__mux2_1 _6289_ (.A0(_3148_),
    .A1(_3288_),
    .S(net213),
    .X(_3289_));
 sky130_fd_sc_hd__o2bb2a_1 _6290_ (.A1_N(_2723_),
    .A2_N(_2986_),
    .B1(_3289_),
    .B2(net186),
    .X(_3290_));
 sky130_fd_sc_hd__a221o_1 _6291_ (.A1(_1502_),
    .A2(net361),
    .B1(net356),
    .B2(_1506_),
    .C1(net363),
    .X(_3291_));
 sky130_fd_sc_hd__o31a_1 _6292_ (.A1(net184),
    .A2(_2989_),
    .A3(_2990_),
    .B1(_3132_),
    .X(_3292_));
 sky130_fd_sc_hd__a22o_1 _6293_ (.A1(_2990_),
    .A2(_3152_),
    .B1(_3291_),
    .B2(_1507_),
    .X(_3293_));
 sky130_fd_sc_hd__or3_1 _6294_ (.A(net222),
    .B(_3290_),
    .C(_3293_),
    .X(_3294_));
 sky130_fd_sc_hd__nand2_1 _6295_ (.A(net2302),
    .B(net222),
    .Y(_3295_));
 sky130_fd_sc_hd__o311a_1 _6296_ (.A1(_3286_),
    .A2(_3292_),
    .A3(_3294_),
    .B1(_3295_),
    .C1(net438),
    .X(_0741_));
 sky130_fd_sc_hd__xnor2_1 _6297_ (.A(_1479_),
    .B(net358),
    .Y(_3296_));
 sky130_fd_sc_hd__and2_1 _6298_ (.A(_1482_),
    .B(_3296_),
    .X(_3297_));
 sky130_fd_sc_hd__nand2_1 _6299_ (.A(_1482_),
    .B(_3296_),
    .Y(_3298_));
 sky130_fd_sc_hd__nor2_1 _6300_ (.A(_1482_),
    .B(_3296_),
    .Y(_3299_));
 sky130_fd_sc_hd__nor2_1 _6301_ (.A(_3297_),
    .B(_3299_),
    .Y(_3300_));
 sky130_fd_sc_hd__a21o_1 _6302_ (.A1(_3279_),
    .A2(_3281_),
    .B1(_3282_),
    .X(_3301_));
 sky130_fd_sc_hd__xnor2_1 _6303_ (.A(_3300_),
    .B(_3301_),
    .Y(_3302_));
 sky130_fd_sc_hd__mux4_1 _6304_ (.A0(_1468_),
    .A1(_1482_),
    .A2(_1447_),
    .A3(_1505_),
    .S0(net199),
    .S1(net191),
    .X(_3303_));
 sky130_fd_sc_hd__or2_1 _6305_ (.A(net202),
    .B(_3303_),
    .X(_3304_));
 sky130_fd_sc_hd__o211a_1 _6306_ (.A1(net206),
    .A2(_3238_),
    .B1(_3304_),
    .C1(net213),
    .X(_3305_));
 sky130_fd_sc_hd__a211o_1 _6307_ (.A1(net209),
    .A2(_3166_),
    .B1(_3305_),
    .C1(net185),
    .X(_3306_));
 sky130_fd_sc_hd__o211a_1 _6308_ (.A1(net189),
    .A2(_3009_),
    .B1(_3306_),
    .C1(_2720_),
    .X(_3307_));
 sky130_fd_sc_hd__nand2_1 _6309_ (.A(net188),
    .B(_3015_),
    .Y(_3308_));
 sky130_fd_sc_hd__a221o_1 _6310_ (.A1(_1483_),
    .A2(net363),
    .B1(net361),
    .B2(_1479_),
    .C1(net222),
    .X(_3309_));
 sky130_fd_sc_hd__nor2_1 _6311_ (.A(net184),
    .B(_2941_),
    .Y(_3310_));
 sky130_fd_sc_hd__a221o_1 _6312_ (.A1(net356),
    .A2(_3300_),
    .B1(_3310_),
    .B2(_2761_),
    .C1(_3309_),
    .X(_3311_));
 sky130_fd_sc_hd__a221o_1 _6313_ (.A1(net317),
    .A2(_3302_),
    .B1(_3308_),
    .B2(_3132_),
    .C1(_3311_),
    .X(_3312_));
 sky130_fd_sc_hd__a21o_1 _6314_ (.A1(net2283),
    .A2(_1482_),
    .B1(net221),
    .X(_3313_));
 sky130_fd_sc_hd__o211a_1 _6315_ (.A1(_3307_),
    .A2(_3312_),
    .B1(net2284),
    .C1(net437),
    .X(_0742_));
 sky130_fd_sc_hd__a21o_1 _6316_ (.A1(_3298_),
    .A2(_3301_),
    .B1(_3299_),
    .X(_3314_));
 sky130_fd_sc_hd__xnor2_1 _6317_ (.A(_1490_),
    .B(net358),
    .Y(_3315_));
 sky130_fd_sc_hd__nor2_1 _6318_ (.A(_1492_),
    .B(_3315_),
    .Y(_3316_));
 sky130_fd_sc_hd__nand2_1 _6319_ (.A(_1492_),
    .B(_3315_),
    .Y(_3317_));
 sky130_fd_sc_hd__nand2b_1 _6320_ (.A_N(_3316_),
    .B(_3317_),
    .Y(_3318_));
 sky130_fd_sc_hd__xnor2_1 _6321_ (.A(_3314_),
    .B(_3318_),
    .Y(_3319_));
 sky130_fd_sc_hd__mux4_1 _6322_ (.A0(_1492_),
    .A1(_1505_),
    .A2(_1482_),
    .A3(_1468_),
    .S0(net196),
    .S1(net191),
    .X(_3320_));
 sky130_fd_sc_hd__mux2_1 _6323_ (.A0(_3254_),
    .A1(_3320_),
    .S(net204),
    .X(_3321_));
 sky130_fd_sc_hd__mux2_1 _6324_ (.A0(_3187_),
    .A1(_3321_),
    .S(net214),
    .X(_3322_));
 sky130_fd_sc_hd__a2bb2o_1 _6325_ (.A1_N(net184),
    .A2_N(_3322_),
    .B1(_3029_),
    .B2(_2723_),
    .X(_3323_));
 sky130_fd_sc_hd__a21oi_1 _6326_ (.A1(net188),
    .A2(_3035_),
    .B1(_3133_),
    .Y(_3324_));
 sky130_fd_sc_hd__nor2_1 _6327_ (.A(net185),
    .B(_3034_),
    .Y(_3325_));
 sky130_fd_sc_hd__a2bb2o_1 _6328_ (.A1_N(_2734_),
    .A2_N(_1493_),
    .B1(_1490_),
    .B2(net361),
    .X(_3326_));
 sky130_fd_sc_hd__o22a_1 _6329_ (.A1(_1490_),
    .A2(_1492_),
    .B1(net363),
    .B2(_3326_),
    .X(_3327_));
 sky130_fd_sc_hd__o21ai_1 _6330_ (.A1(_2731_),
    .A2(_3319_),
    .B1(_3323_),
    .Y(_3328_));
 sky130_fd_sc_hd__or4_1 _6331_ (.A(net222),
    .B(_3325_),
    .C(_3327_),
    .D(_3328_),
    .X(_3329_));
 sky130_fd_sc_hd__o221a_1 _6332_ (.A1(_1493_),
    .A2(net221),
    .B1(_3324_),
    .B2(_3329_),
    .C1(net437),
    .X(_0743_));
 sky130_fd_sc_hd__xnor2_1 _6333_ (.A(_1514_),
    .B(net358),
    .Y(_3330_));
 sky130_fd_sc_hd__nor2_1 _6334_ (.A(_1516_),
    .B(_3330_),
    .Y(_3331_));
 sky130_fd_sc_hd__nand2_1 _6335_ (.A(_1516_),
    .B(_3330_),
    .Y(_3332_));
 sky130_fd_sc_hd__and2b_1 _6336_ (.A_N(_3331_),
    .B(_3332_),
    .X(_3333_));
 sky130_fd_sc_hd__a21o_1 _6337_ (.A1(_3314_),
    .A2(_3317_),
    .B1(_3316_),
    .X(_3334_));
 sky130_fd_sc_hd__nand2_1 _6338_ (.A(_3333_),
    .B(_3334_),
    .Y(_3335_));
 sky130_fd_sc_hd__or2_1 _6339_ (.A(_3333_),
    .B(_3334_),
    .X(_3336_));
 sky130_fd_sc_hd__a21oi_1 _6340_ (.A1(_3335_),
    .A2(_3336_),
    .B1(_2731_),
    .Y(_3337_));
 sky130_fd_sc_hd__mux4_1 _6341_ (.A0(_1482_),
    .A1(_1505_),
    .A2(_1516_),
    .A3(_1492_),
    .S0(net191),
    .S1(net199),
    .X(_3338_));
 sky130_fd_sc_hd__mux2_1 _6342_ (.A0(_3273_),
    .A1(_3338_),
    .S(net204),
    .X(_3339_));
 sky130_fd_sc_hd__mux2_1 _6343_ (.A0(_3200_),
    .A1(_3339_),
    .S(net212),
    .X(_3340_));
 sky130_fd_sc_hd__o2bb2a_1 _6344_ (.A1_N(_2723_),
    .A2_N(_3049_),
    .B1(_3340_),
    .B2(net184),
    .X(_3341_));
 sky130_fd_sc_hd__nand2_1 _6345_ (.A(net188),
    .B(_3054_),
    .Y(_3342_));
 sky130_fd_sc_hd__a21o_1 _6346_ (.A1(_1514_),
    .A2(net361),
    .B1(net363),
    .X(_3343_));
 sky130_fd_sc_hd__o21a_1 _6347_ (.A1(_1514_),
    .A2(_1516_),
    .B1(_3343_),
    .X(_3344_));
 sky130_fd_sc_hd__a211o_1 _6348_ (.A1(net356),
    .A2(_3333_),
    .B1(_3344_),
    .C1(net222),
    .X(_3345_));
 sky130_fd_sc_hd__a221o_1 _6349_ (.A1(_2839_),
    .A2(_3310_),
    .B1(_3342_),
    .B2(_3132_),
    .C1(_3345_),
    .X(_3346_));
 sky130_fd_sc_hd__a21o_1 _6350_ (.A1(_1514_),
    .A2(net2331),
    .B1(net221),
    .X(_3347_));
 sky130_fd_sc_hd__o311a_1 _6351_ (.A1(_3337_),
    .A2(_3341_),
    .A3(_3346_),
    .B1(_3347_),
    .C1(net437),
    .X(_0744_));
 sky130_fd_sc_hd__a21o_1 _6352_ (.A1(_3332_),
    .A2(_3334_),
    .B1(_3331_),
    .X(_3348_));
 sky130_fd_sc_hd__xnor2_1 _6353_ (.A(_1347_),
    .B(net358),
    .Y(_3349_));
 sky130_fd_sc_hd__nor2_1 _6354_ (.A(_1350_),
    .B(_3349_),
    .Y(_3350_));
 sky130_fd_sc_hd__nand2_1 _6355_ (.A(_1350_),
    .B(_3349_),
    .Y(_3351_));
 sky130_fd_sc_hd__nand2b_1 _6356_ (.A_N(_3350_),
    .B(_3351_),
    .Y(_3352_));
 sky130_fd_sc_hd__xnor2_1 _6357_ (.A(_3348_),
    .B(_3352_),
    .Y(_3353_));
 sky130_fd_sc_hd__mux4_1 _6358_ (.A0(_1350_),
    .A1(_1492_),
    .A2(_1516_),
    .A3(_1482_),
    .S0(net196),
    .S1(net191),
    .X(_3354_));
 sky130_fd_sc_hd__mux2_1 _6359_ (.A0(_3287_),
    .A1(_3354_),
    .S(net206),
    .X(_3355_));
 sky130_fd_sc_hd__mux2_1 _6360_ (.A0(_3218_),
    .A1(_3355_),
    .S(net213),
    .X(_3356_));
 sky130_fd_sc_hd__nor2_1 _6361_ (.A(net186),
    .B(_3356_),
    .Y(_3357_));
 sky130_fd_sc_hd__a211o_1 _6362_ (.A1(net186),
    .A2(_3070_),
    .B1(_3357_),
    .C1(_2721_),
    .X(_3358_));
 sky130_fd_sc_hd__a21o_1 _6363_ (.A1(net188),
    .A2(_3075_),
    .B1(_3133_),
    .X(_3359_));
 sky130_fd_sc_hd__a221o_1 _6364_ (.A1(_1347_),
    .A2(net361),
    .B1(net356),
    .B2(_1351_),
    .C1(net363),
    .X(_3360_));
 sky130_fd_sc_hd__a21o_1 _6365_ (.A1(_1352_),
    .A2(_3360_),
    .B1(net222),
    .X(_3361_));
 sky130_fd_sc_hd__a21oi_1 _6366_ (.A1(_2873_),
    .A2(_3310_),
    .B1(_3361_),
    .Y(_3362_));
 sky130_fd_sc_hd__o2111a_1 _6367_ (.A1(_2731_),
    .A2(_3353_),
    .B1(_3358_),
    .C1(_3359_),
    .D1(_3362_),
    .X(_3363_));
 sky130_fd_sc_hd__a211oi_1 _6368_ (.A1(net2271),
    .A2(net222),
    .B1(_3363_),
    .C1(net466),
    .Y(_0745_));
 sky130_fd_sc_hd__xnor2_1 _6369_ (.A(_1370_),
    .B(net358),
    .Y(_3364_));
 sky130_fd_sc_hd__nor2_1 _6370_ (.A(_1373_),
    .B(_3364_),
    .Y(_3365_));
 sky130_fd_sc_hd__nand2_1 _6371_ (.A(_1373_),
    .B(_3364_),
    .Y(_3366_));
 sky130_fd_sc_hd__and2b_1 _6372_ (.A_N(_3365_),
    .B(_3366_),
    .X(_3367_));
 sky130_fd_sc_hd__a21o_1 _6373_ (.A1(_3348_),
    .A2(_3351_),
    .B1(_3350_),
    .X(_3368_));
 sky130_fd_sc_hd__xor2_1 _6374_ (.A(_3367_),
    .B(_3368_),
    .X(_3369_));
 sky130_fd_sc_hd__nor2_1 _6375_ (.A(_2731_),
    .B(_3369_),
    .Y(_3370_));
 sky130_fd_sc_hd__mux4_1 _6376_ (.A0(_1373_),
    .A1(_1516_),
    .A2(_1350_),
    .A3(_1492_),
    .S0(net196),
    .S1(net191),
    .X(_3371_));
 sky130_fd_sc_hd__mux2_1 _6377_ (.A0(_3303_),
    .A1(_3371_),
    .S(net204),
    .X(_3372_));
 sky130_fd_sc_hd__mux2_1 _6378_ (.A0(_3239_),
    .A1(_3372_),
    .S(net213),
    .X(_3373_));
 sky130_fd_sc_hd__o2bb2a_1 _6379_ (.A1_N(_2723_),
    .A2_N(_3092_),
    .B1(_3373_),
    .B2(net185),
    .X(_3374_));
 sky130_fd_sc_hd__a21oi_1 _6380_ (.A1(net188),
    .A2(_3097_),
    .B1(_3133_),
    .Y(_3375_));
 sky130_fd_sc_hd__a221o_1 _6381_ (.A1(_1374_),
    .A2(net363),
    .B1(net361),
    .B2(_1370_),
    .C1(net222),
    .X(_3376_));
 sky130_fd_sc_hd__a32o_1 _6382_ (.A1(net188),
    .A2(_2898_),
    .A3(_2940_),
    .B1(_3367_),
    .B2(net356),
    .X(_3377_));
 sky130_fd_sc_hd__or4_1 _6383_ (.A(_3374_),
    .B(_3375_),
    .C(_3376_),
    .D(_3377_),
    .X(_3378_));
 sky130_fd_sc_hd__a21o_1 _6384_ (.A1(_1370_),
    .A2(_1373_),
    .B1(net221),
    .X(_3379_));
 sky130_fd_sc_hd__o211a_1 _6385_ (.A1(_3370_),
    .A2(_3378_),
    .B1(net2261),
    .C1(net437),
    .X(_0746_));
 sky130_fd_sc_hd__a21o_1 _6386_ (.A1(_3366_),
    .A2(_3368_),
    .B1(_3365_),
    .X(_3380_));
 sky130_fd_sc_hd__xnor2_1 _6387_ (.A(_1358_),
    .B(_2729_),
    .Y(_3381_));
 sky130_fd_sc_hd__inv_2 _6388_ (.A(_3381_),
    .Y(_3382_));
 sky130_fd_sc_hd__nor2_1 _6389_ (.A(_1360_),
    .B(_3382_),
    .Y(_3383_));
 sky130_fd_sc_hd__nand2_1 _6390_ (.A(_1360_),
    .B(_3382_),
    .Y(_3384_));
 sky130_fd_sc_hd__nand2b_1 _6391_ (.A_N(_3383_),
    .B(_3384_),
    .Y(_3385_));
 sky130_fd_sc_hd__xnor2_1 _6392_ (.A(_3380_),
    .B(_3385_),
    .Y(_3386_));
 sky130_fd_sc_hd__mux4_1 _6393_ (.A0(_1350_),
    .A1(_1360_),
    .A2(_1516_),
    .A3(_1373_),
    .S0(net199),
    .S1(net195),
    .X(_3387_));
 sky130_fd_sc_hd__mux2_1 _6394_ (.A0(_3320_),
    .A1(_3387_),
    .S(net204),
    .X(_3388_));
 sky130_fd_sc_hd__mux2_1 _6395_ (.A0(_3255_),
    .A1(_3388_),
    .S(net214),
    .X(_3389_));
 sky130_fd_sc_hd__a2bb2o_1 _6396_ (.A1_N(net184),
    .A2_N(_3389_),
    .B1(_3111_),
    .B2(_2723_),
    .X(_3390_));
 sky130_fd_sc_hd__a21oi_1 _6397_ (.A1(net188),
    .A2(_3116_),
    .B1(_3133_),
    .Y(_3391_));
 sky130_fd_sc_hd__a221o_1 _6398_ (.A1(_1358_),
    .A2(net361),
    .B1(net356),
    .B2(_1361_),
    .C1(net363),
    .X(_3392_));
 sky130_fd_sc_hd__o21a_1 _6399_ (.A1(_1358_),
    .A2(_1360_),
    .B1(_3392_),
    .X(_3393_));
 sky130_fd_sc_hd__a2111oi_1 _6400_ (.A1(_2942_),
    .A2(_3310_),
    .B1(_3391_),
    .C1(_3393_),
    .D1(net222),
    .Y(_3394_));
 sky130_fd_sc_hd__o211a_1 _6401_ (.A1(_2731_),
    .A2(_3386_),
    .B1(_3390_),
    .C1(_3394_),
    .X(_3395_));
 sky130_fd_sc_hd__a211oi_4 _6402_ (.A1(_1361_),
    .A2(net222),
    .B1(_3395_),
    .C1(net466),
    .Y(_0747_));
 sky130_fd_sc_hd__a21oi_1 _6403_ (.A1(_3380_),
    .A2(_3384_),
    .B1(_3383_),
    .Y(_3396_));
 sky130_fd_sc_hd__and2_1 _6404_ (.A(_1339_),
    .B(net358),
    .X(_3397_));
 sky130_fd_sc_hd__nor2_1 _6405_ (.A(_1339_),
    .B(net358),
    .Y(_3398_));
 sky130_fd_sc_hd__nor2_1 _6406_ (.A(_3397_),
    .B(_3398_),
    .Y(_3399_));
 sky130_fd_sc_hd__a211o_1 _6407_ (.A1(_3380_),
    .A2(_3384_),
    .B1(_3399_),
    .C1(_3383_),
    .X(_3400_));
 sky130_fd_sc_hd__o311a_1 _6408_ (.A1(_3396_),
    .A2(_3397_),
    .A3(_3398_),
    .B1(_3400_),
    .C1(net317),
    .X(_3401_));
 sky130_fd_sc_hd__mux4_1 _6409_ (.A0(_1337_),
    .A1(_1360_),
    .A2(_1373_),
    .A3(_1350_),
    .S0(net191),
    .S1(net197),
    .X(_3402_));
 sky130_fd_sc_hd__or2_1 _6410_ (.A(net201),
    .B(_3402_),
    .X(_3403_));
 sky130_fd_sc_hd__o211a_1 _6411_ (.A1(net204),
    .A2(_3338_),
    .B1(_3403_),
    .C1(net212),
    .X(_3404_));
 sky130_fd_sc_hd__a211o_1 _6412_ (.A1(net208),
    .A2(_3274_),
    .B1(_3404_),
    .C1(net185),
    .X(_3405_));
 sky130_fd_sc_hd__o211a_1 _6413_ (.A1(net189),
    .A2(_3129_),
    .B1(_3405_),
    .C1(_2720_),
    .X(_3406_));
 sky130_fd_sc_hd__o21a_1 _6414_ (.A1(_1321_),
    .A2(_1337_),
    .B1(net363),
    .X(_3407_));
 sky130_fd_sc_hd__a221o_1 _6415_ (.A1(_1337_),
    .A2(_2686_),
    .B1(net361),
    .B2(_1321_),
    .C1(net222),
    .X(_3408_));
 sky130_fd_sc_hd__a211o_1 _6416_ (.A1(_1339_),
    .A2(net356),
    .B1(_3407_),
    .C1(_3408_),
    .X(_3409_));
 sky130_fd_sc_hd__a31o_1 _6417_ (.A1(net211),
    .A2(_2970_),
    .A3(_3152_),
    .B1(_3409_),
    .X(_3410_));
 sky130_fd_sc_hd__a21o_1 _6418_ (.A1(_1321_),
    .A2(_1337_),
    .B1(net221),
    .X(_3411_));
 sky130_fd_sc_hd__o311a_1 _6419_ (.A1(_3401_),
    .A2(_3406_),
    .A3(_3410_),
    .B1(net2278),
    .C1(net437),
    .X(_0748_));
 sky130_fd_sc_hd__and2_1 _6420_ (.A(net1987),
    .B(net443),
    .X(_0749_));
 sky130_fd_sc_hd__and2_1 _6421_ (.A(net610),
    .B(net443),
    .X(_0750_));
 sky130_fd_sc_hd__and2_1 _6422_ (.A(net452),
    .B(net739),
    .X(_0751_));
 sky130_fd_sc_hd__and2_1 _6423_ (.A(net445),
    .B(_1566_),
    .X(_0752_));
 sky130_fd_sc_hd__o31a_2 _6424_ (.A1(_1549_),
    .A2(_1550_),
    .A3(_1551_),
    .B1(net443),
    .X(_0753_));
 sky130_fd_sc_hd__and2_1 _6425_ (.A(net444),
    .B(_1537_),
    .X(_0754_));
 sky130_fd_sc_hd__nor2_1 _6426_ (.A(net471),
    .B(_1525_),
    .Y(_0755_));
 sky130_fd_sc_hd__and2_1 _6427_ (.A(net459),
    .B(_1586_),
    .X(_0756_));
 sky130_fd_sc_hd__o31a_1 _6428_ (.A1(_1609_),
    .A2(_1610_),
    .A3(_1611_),
    .B1(net451),
    .X(_0757_));
 sky130_fd_sc_hd__and2_1 _6429_ (.A(net458),
    .B(_1598_),
    .X(_0758_));
 sky130_fd_sc_hd__and2_1 _6430_ (.A(net447),
    .B(net2251),
    .X(_0759_));
 sky130_fd_sc_hd__nor2_1 _6431_ (.A(net466),
    .B(_1646_),
    .Y(_0760_));
 sky130_fd_sc_hd__and2_1 _6432_ (.A(net451),
    .B(_1626_),
    .X(_0761_));
 sky130_fd_sc_hd__and2_1 _6433_ (.A(net456),
    .B(_1635_),
    .X(_0762_));
 sky130_fd_sc_hd__and2_1 _6434_ (.A(net438),
    .B(_1657_),
    .X(_0763_));
 sky130_fd_sc_hd__nor2_1 _6435_ (.A(net468),
    .B(_1692_),
    .Y(_0764_));
 sky130_fd_sc_hd__and2_1 _6436_ (.A(net440),
    .B(_1669_),
    .X(_0765_));
 sky130_fd_sc_hd__and2_1 _6437_ (.A(net444),
    .B(_1681_),
    .X(_0766_));
 sky130_fd_sc_hd__and2_1 _6438_ (.A(net437),
    .B(_1704_),
    .X(_0767_));
 sky130_fd_sc_hd__nor2_2 _6439_ (.A(net468),
    .B(_1409_),
    .Y(_0768_));
 sky130_fd_sc_hd__a31oi_2 _6440_ (.A1(_1383_),
    .A2(_1384_),
    .A3(_1385_),
    .B1(net467),
    .Y(_0769_));
 sky130_fd_sc_hd__and2_1 _6441_ (.A(net458),
    .B(_1422_),
    .X(_0770_));
 sky130_fd_sc_hd__and2_1 _6442_ (.A(net444),
    .B(_1398_),
    .X(_0771_));
 sky130_fd_sc_hd__nor2_1 _6443_ (.A(net467),
    .B(_1454_),
    .Y(_0772_));
 sky130_fd_sc_hd__and2_1 _6444_ (.A(net441),
    .B(_1434_),
    .X(_0773_));
 sky130_fd_sc_hd__and2_2 _6445_ (.A(net453),
    .B(_1444_),
    .X(_0774_));
 sky130_fd_sc_hd__and2_1 _6446_ (.A(net441),
    .B(_1465_),
    .X(_0775_));
 sky130_fd_sc_hd__nor2_1 _6447_ (.A(net471),
    .B(_1500_),
    .Y(_0776_));
 sky130_fd_sc_hd__nor2_1 _6448_ (.A(net467),
    .B(_1477_),
    .Y(_0777_));
 sky130_fd_sc_hd__and2_1 _6449_ (.A(net437),
    .B(_1489_),
    .X(_0778_));
 sky130_fd_sc_hd__nor2_1 _6450_ (.A(net469),
    .B(_1512_),
    .Y(_0779_));
 sky130_fd_sc_hd__nor2_1 _6451_ (.A(net466),
    .B(_1345_),
    .Y(_0780_));
 sky130_fd_sc_hd__nor2_1 _6452_ (.A(net466),
    .B(net2222),
    .Y(_0781_));
 sky130_fd_sc_hd__and2_1 _6453_ (.A(net453),
    .B(_1357_),
    .X(_0782_));
 sky130_fd_sc_hd__nor2_1 _6454_ (.A(net464),
    .B(_1319_),
    .Y(_0783_));
 sky130_fd_sc_hd__and2_1 _6455_ (.A(net443),
    .B(net2037),
    .X(_0784_));
 sky130_fd_sc_hd__and2_1 _6456_ (.A(net459),
    .B(net596),
    .X(_0785_));
 sky130_fd_sc_hd__and2_1 _6457_ (.A(net459),
    .B(net748),
    .X(_0786_));
 sky130_fd_sc_hd__and2_1 _6458_ (.A(net437),
    .B(net2105),
    .X(_0787_));
 sky130_fd_sc_hd__and2_1 _6459_ (.A(net2109),
    .B(net455),
    .X(_0788_));
 sky130_fd_sc_hd__mux2_1 _6460_ (.A0(net2062),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .S(net472),
    .X(_0789_));
 sky130_fd_sc_hd__mux2_1 _6461_ (.A0(net2038),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .S(net472),
    .X(_0790_));
 sky130_fd_sc_hd__mux2_1 _6462_ (.A0(net1982),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .S(net472),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _6463_ (.A0(net1985),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .S(net472),
    .X(_0792_));
 sky130_fd_sc_hd__and2_1 _6464_ (.A(net438),
    .B(net770),
    .X(_0793_));
 sky130_fd_sc_hd__and2_1 _6465_ (.A(net451),
    .B(net586),
    .X(_0794_));
 sky130_fd_sc_hd__and2_1 _6466_ (.A(net451),
    .B(net626),
    .X(_0795_));
 sky130_fd_sc_hd__and2_1 _6467_ (.A(net451),
    .B(net584),
    .X(_0796_));
 sky130_fd_sc_hd__and2_1 _6468_ (.A(net449),
    .B(net689),
    .X(_0797_));
 sky130_fd_sc_hd__and2_1 _6469_ (.A(net457),
    .B(net733),
    .X(_0798_));
 sky130_fd_sc_hd__and2_1 _6470_ (.A(net457),
    .B(net709),
    .X(_0799_));
 sky130_fd_sc_hd__and2_1 _6471_ (.A(net457),
    .B(net598),
    .X(_0800_));
 sky130_fd_sc_hd__and2_1 _6472_ (.A(net449),
    .B(net624),
    .X(_0801_));
 sky130_fd_sc_hd__and2_1 _6473_ (.A(net443),
    .B(net652),
    .X(_0802_));
 sky130_fd_sc_hd__and2_1 _6474_ (.A(net457),
    .B(net750),
    .X(_0803_));
 sky130_fd_sc_hd__and2_1 _6475_ (.A(net449),
    .B(net604),
    .X(_0804_));
 sky130_fd_sc_hd__and2_1 _6476_ (.A(net449),
    .B(net618),
    .X(_0805_));
 sky130_fd_sc_hd__and2_1 _6477_ (.A(net449),
    .B(net574),
    .X(_0806_));
 sky130_fd_sc_hd__and2_1 _6478_ (.A(net453),
    .B(net662),
    .X(_0807_));
 sky130_fd_sc_hd__and2_1 _6479_ (.A(net450),
    .B(net727),
    .X(_0808_));
 sky130_fd_sc_hd__and2_1 _6480_ (.A(net455),
    .B(net564),
    .X(_0809_));
 sky130_fd_sc_hd__and2_1 _6481_ (.A(net447),
    .B(net705),
    .X(_0810_));
 sky130_fd_sc_hd__and2_1 _6482_ (.A(net441),
    .B(net654),
    .X(_0811_));
 sky130_fd_sc_hd__and2_1 _6483_ (.A(net442),
    .B(net628),
    .X(_0812_));
 sky130_fd_sc_hd__and2_1 _6484_ (.A(net441),
    .B(net681),
    .X(_0813_));
 sky130_fd_sc_hd__and2_1 _6485_ (.A(net442),
    .B(net701),
    .X(_0814_));
 sky130_fd_sc_hd__and2_1 _6486_ (.A(net441),
    .B(net723),
    .X(_0815_));
 sky130_fd_sc_hd__and2_1 _6487_ (.A(net440),
    .B(net699),
    .X(_0816_));
 sky130_fd_sc_hd__and2_1 _6488_ (.A(net440),
    .B(net683),
    .X(_0817_));
 sky130_fd_sc_hd__and2_1 _6489_ (.A(net440),
    .B(net592),
    .X(_0818_));
 sky130_fd_sc_hd__and2_1 _6490_ (.A(net437),
    .B(net768),
    .X(_0819_));
 sky130_fd_sc_hd__and2_1 _6491_ (.A(net439),
    .B(net1476),
    .X(_0820_));
 sky130_fd_sc_hd__and2_1 _6492_ (.A(net439),
    .B(net766),
    .X(_0821_));
 sky130_fd_sc_hd__and2_1 _6493_ (.A(net440),
    .B(net594),
    .X(_0822_));
 sky130_fd_sc_hd__and2_1 _6494_ (.A(net453),
    .B(net568),
    .X(_0823_));
 sky130_fd_sc_hd__and2_1 _6495_ (.A(net444),
    .B(net550),
    .X(_0824_));
 sky130_fd_sc_hd__and2_1 _6496_ (.A(net438),
    .B(net746),
    .X(_0825_));
 sky130_fd_sc_hd__and2_1 _6497_ (.A(net452),
    .B(net703),
    .X(_0826_));
 sky130_fd_sc_hd__and2_1 _6498_ (.A(net457),
    .B(net622),
    .X(_0827_));
 sky130_fd_sc_hd__and2_1 _6499_ (.A(net451),
    .B(net675),
    .X(_0828_));
 sky130_fd_sc_hd__and2_1 _6500_ (.A(net450),
    .B(net616),
    .X(_0829_));
 sky130_fd_sc_hd__and2_1 _6501_ (.A(net458),
    .B(net721),
    .X(_0830_));
 sky130_fd_sc_hd__and2_1 _6502_ (.A(net457),
    .B(net612),
    .X(_0831_));
 sky130_fd_sc_hd__and2_1 _6503_ (.A(net457),
    .B(net673),
    .X(_0832_));
 sky130_fd_sc_hd__and2_1 _6504_ (.A(net450),
    .B(net572),
    .X(_0833_));
 sky130_fd_sc_hd__and2_1 _6505_ (.A(net449),
    .B(net687),
    .X(_0834_));
 sky130_fd_sc_hd__and2_1 _6506_ (.A(net457),
    .B(net606),
    .X(_0835_));
 sky130_fd_sc_hd__and2_1 _6507_ (.A(net449),
    .B(net644),
    .X(_0836_));
 sky130_fd_sc_hd__and2_1 _6508_ (.A(net449),
    .B(net664),
    .X(_0837_));
 sky130_fd_sc_hd__and2_1 _6509_ (.A(net449),
    .B(net668),
    .X(_0838_));
 sky130_fd_sc_hd__and2_1 _6510_ (.A(net453),
    .B(net630),
    .X(_0839_));
 sky130_fd_sc_hd__and2_1 _6511_ (.A(net450),
    .B(net685),
    .X(_0840_));
 sky130_fd_sc_hd__and2_1 _6512_ (.A(net455),
    .B(net758),
    .X(_0841_));
 sky130_fd_sc_hd__and2_1 _6513_ (.A(net443),
    .B(net693),
    .X(_0842_));
 sky130_fd_sc_hd__and2_1 _6514_ (.A(net441),
    .B(net562),
    .X(_0843_));
 sky130_fd_sc_hd__and2_1 _6515_ (.A(net442),
    .B(net632),
    .X(_0844_));
 sky130_fd_sc_hd__and2_1 _6516_ (.A(net441),
    .B(net558),
    .X(_0845_));
 sky130_fd_sc_hd__and2_1 _6517_ (.A(net442),
    .B(net719),
    .X(_0846_));
 sky130_fd_sc_hd__and2_1 _6518_ (.A(net441),
    .B(net640),
    .X(_0847_));
 sky130_fd_sc_hd__and2_1 _6519_ (.A(net440),
    .B(net620),
    .X(_0848_));
 sky130_fd_sc_hd__and2_1 _6520_ (.A(net439),
    .B(net638),
    .X(_0849_));
 sky130_fd_sc_hd__and2_1 _6521_ (.A(net440),
    .B(net578),
    .X(_0850_));
 sky130_fd_sc_hd__and2_1 _6522_ (.A(net439),
    .B(net560),
    .X(_0851_));
 sky130_fd_sc_hd__and2_1 _6523_ (.A(net439),
    .B(net590),
    .X(_0852_));
 sky130_fd_sc_hd__and2_1 _6524_ (.A(net439),
    .B(net642),
    .X(_0853_));
 sky130_fd_sc_hd__and2_1 _6525_ (.A(net439),
    .B(net570),
    .X(_0854_));
 sky130_fd_sc_hd__and2_1 _6526_ (.A(net2007),
    .B(net453),
    .X(_0855_));
 sky130_fd_sc_hd__nor2_1 _6527_ (.A(_1290_),
    .B(net467),
    .Y(_0856_));
 sky130_fd_sc_hd__and2_1 _6528_ (.A(net860),
    .B(net437),
    .X(_0857_));
 sky130_fd_sc_hd__and2_1 _6529_ (.A(net1984),
    .B(net451),
    .X(_0858_));
 sky130_fd_sc_hd__and2_1 _6530_ (.A(net1928),
    .B(net457),
    .X(_0859_));
 sky130_fd_sc_hd__and2_1 _6531_ (.A(net2152),
    .B(net452),
    .X(_0860_));
 sky130_fd_sc_hd__and2_1 _6532_ (.A(net2067),
    .B(net450),
    .X(_0861_));
 sky130_fd_sc_hd__and2_1 _6533_ (.A(net2034),
    .B(net451),
    .X(_0862_));
 sky130_fd_sc_hd__and2_1 _6534_ (.A(net2008),
    .B(net452),
    .X(_0863_));
 sky130_fd_sc_hd__and2_1 _6535_ (.A(net2104),
    .B(net458),
    .X(_0864_));
 sky130_fd_sc_hd__and2_1 _6536_ (.A(net962),
    .B(net450),
    .X(_0865_));
 sky130_fd_sc_hd__and2_1 _6537_ (.A(net778),
    .B(net443),
    .X(_0866_));
 sky130_fd_sc_hd__and2_1 _6538_ (.A(net2130),
    .B(net457),
    .X(_0867_));
 sky130_fd_sc_hd__and2_1 _6539_ (.A(net1855),
    .B(net453),
    .X(_0868_));
 sky130_fd_sc_hd__and2_1 _6540_ (.A(net2147),
    .B(net450),
    .X(_0869_));
 sky130_fd_sc_hd__and2_1 _6541_ (.A(net2129),
    .B(net451),
    .X(_0870_));
 sky130_fd_sc_hd__and2_1 _6542_ (.A(net2047),
    .B(net454),
    .X(_0871_));
 sky130_fd_sc_hd__and2_1 _6543_ (.A(net898),
    .B(net443),
    .X(_0872_));
 sky130_fd_sc_hd__and2_1 _6544_ (.A(net1977),
    .B(net455),
    .X(_0873_));
 sky130_fd_sc_hd__and2_1 _6545_ (.A(net2168),
    .B(net443),
    .X(_0874_));
 sky130_fd_sc_hd__and2_1 _6546_ (.A(net2080),
    .B(net441),
    .X(_0875_));
 sky130_fd_sc_hd__and2_1 _6547_ (.A(net2005),
    .B(net442),
    .X(_0876_));
 sky130_fd_sc_hd__and2_1 _6548_ (.A(net2185),
    .B(net441),
    .X(_0877_));
 sky130_fd_sc_hd__and2_1 _6549_ (.A(net2016),
    .B(net442),
    .X(_0878_));
 sky130_fd_sc_hd__and2_1 _6550_ (.A(net2159),
    .B(net441),
    .X(_0879_));
 sky130_fd_sc_hd__and2_1 _6551_ (.A(net2006),
    .B(net442),
    .X(_0880_));
 sky130_fd_sc_hd__and2_1 _6552_ (.A(net2143),
    .B(net442),
    .X(_0881_));
 sky130_fd_sc_hd__and2_1 _6553_ (.A(net2178),
    .B(net439),
    .X(_0882_));
 sky130_fd_sc_hd__and2_1 _6554_ (.A(net1996),
    .B(net437),
    .X(_0883_));
 sky130_fd_sc_hd__and2_1 _6555_ (.A(net2198),
    .B(net439),
    .X(_0884_));
 sky130_fd_sc_hd__and2_1 _6556_ (.A(net670),
    .B(net453),
    .X(_0885_));
 sky130_fd_sc_hd__and2_1 _6557_ (.A(net2158),
    .B(net440),
    .X(_0886_));
 sky130_fd_sc_hd__and3_2 _6558_ (.A(net1698),
    .B(net178),
    .C(net280),
    .X(_0887_));
 sky130_fd_sc_hd__and3_1 _6559_ (.A(net1998),
    .B(net180),
    .C(net289),
    .X(_0888_));
 sky130_fd_sc_hd__and3_1 _6560_ (.A(net1990),
    .B(net2232),
    .C(net277),
    .X(_0889_));
 sky130_fd_sc_hd__nor4_2 _6561_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2614_),
    .D(_2637_),
    .Y(_3412_));
 sky130_fd_sc_hd__inv_2 _6562_ (.A(_3412_),
    .Y(_3413_));
 sky130_fd_sc_hd__nor2_2 _6563_ (.A(net471),
    .B(net315),
    .Y(_3414_));
 sky130_fd_sc_hd__or2_1 _6564_ (.A(net471),
    .B(net314),
    .X(_3415_));
 sky130_fd_sc_hd__o22a_1 _6565_ (.A1(net329),
    .A2(_3413_),
    .B1(_3415_),
    .B2(net810),
    .X(_0890_));
 sky130_fd_sc_hd__o22a_1 _6566_ (.A1(net330),
    .A2(_3413_),
    .B1(_3415_),
    .B2(net873),
    .X(_0891_));
 sky130_fd_sc_hd__a22o_1 _6567_ (.A1(net331),
    .A2(net314),
    .B1(net258),
    .B2(net977),
    .X(_0892_));
 sky130_fd_sc_hd__a22o_1 _6568_ (.A1(net332),
    .A2(net314),
    .B1(net257),
    .B2(net1147),
    .X(_0893_));
 sky130_fd_sc_hd__a22o_1 _6569_ (.A1(net327),
    .A2(net314),
    .B1(net258),
    .B2(net1275),
    .X(_0894_));
 sky130_fd_sc_hd__a22o_1 _6570_ (.A1(_1608_),
    .A2(net314),
    .B1(net258),
    .B2(net1556),
    .X(_0895_));
 sky130_fd_sc_hd__a22o_1 _6571_ (.A1(net326),
    .A2(net314),
    .B1(net258),
    .B2(net1197),
    .X(_0896_));
 sky130_fd_sc_hd__a22o_1 _6572_ (.A1(net328),
    .A2(net314),
    .B1(net257),
    .B2(net1722),
    .X(_0897_));
 sky130_fd_sc_hd__a22o_1 _6573_ (.A1(net323),
    .A2(net314),
    .B1(net258),
    .B2(net1139),
    .X(_0898_));
 sky130_fd_sc_hd__a22o_1 _6574_ (.A1(net325),
    .A2(net316),
    .B1(net258),
    .B2(net987),
    .X(_0899_));
 sky130_fd_sc_hd__a22o_1 _6575_ (.A1(net324),
    .A2(net314),
    .B1(net258),
    .B2(net1051),
    .X(_0900_));
 sky130_fd_sc_hd__a22o_1 _6576_ (.A1(net322),
    .A2(net315),
    .B1(net257),
    .B2(net1123),
    .X(_0901_));
 sky130_fd_sc_hd__a22o_1 _6577_ (.A1(net319),
    .A2(net314),
    .B1(net258),
    .B2(net1321),
    .X(_0902_));
 sky130_fd_sc_hd__a22o_1 _6578_ (.A1(net321),
    .A2(net315),
    .B1(net257),
    .B2(net1149),
    .X(_0903_));
 sky130_fd_sc_hd__a22o_1 _6579_ (.A1(net320),
    .A2(net314),
    .B1(net258),
    .B2(net1213),
    .X(_0904_));
 sky130_fd_sc_hd__a22o_1 _6580_ (.A1(net318),
    .A2(net314),
    .B1(net258),
    .B2(net1293),
    .X(_0905_));
 sky130_fd_sc_hd__a22o_1 _6581_ (.A1(net342),
    .A2(net315),
    .B1(net257),
    .B2(net1181),
    .X(_0906_));
 sky130_fd_sc_hd__a22o_1 _6582_ (.A1(_1382_),
    .A2(net315),
    .B1(net257),
    .B2(net905),
    .X(_0907_));
 sky130_fd_sc_hd__a22o_1 _6583_ (.A1(net341),
    .A2(net314),
    .B1(net258),
    .B2(net1145),
    .X(_0908_));
 sky130_fd_sc_hd__a22o_1 _6584_ (.A1(net343),
    .A2(net315),
    .B1(net257),
    .B2(net1067),
    .X(_0909_));
 sky130_fd_sc_hd__a22o_1 _6585_ (.A1(net338),
    .A2(net315),
    .B1(net257),
    .B2(net1313),
    .X(_0910_));
 sky130_fd_sc_hd__a22o_1 _6586_ (.A1(net340),
    .A2(net315),
    .B1(net257),
    .B2(net1245),
    .X(_0911_));
 sky130_fd_sc_hd__a22o_1 _6587_ (.A1(net339),
    .A2(net314),
    .B1(net258),
    .B2(net1413),
    .X(_0912_));
 sky130_fd_sc_hd__a22o_1 _6588_ (.A1(net337),
    .A2(net315),
    .B1(net257),
    .B2(net1726),
    .X(_0913_));
 sky130_fd_sc_hd__a22o_1 _6589_ (.A1(net334),
    .A2(net314),
    .B1(net258),
    .B2(net1750),
    .X(_0914_));
 sky130_fd_sc_hd__a22o_1 _6590_ (.A1(net336),
    .A2(net315),
    .B1(net257),
    .B2(net1189),
    .X(_0915_));
 sky130_fd_sc_hd__a22o_1 _6591_ (.A1(net335),
    .A2(net315),
    .B1(net257),
    .B2(net1522),
    .X(_0916_));
 sky130_fd_sc_hd__a22o_1 _6592_ (.A1(net333),
    .A2(net315),
    .B1(net257),
    .B2(net899),
    .X(_0917_));
 sky130_fd_sc_hd__a22o_1 _6593_ (.A1(net346),
    .A2(net315),
    .B1(net257),
    .B2(net1183),
    .X(_0918_));
 sky130_fd_sc_hd__a22o_1 _6594_ (.A1(net344),
    .A2(net315),
    .B1(net257),
    .B2(net1251),
    .X(_0919_));
 sky130_fd_sc_hd__a22o_1 _6595_ (.A1(net345),
    .A2(net314),
    .B1(net258),
    .B2(net1339),
    .X(_0920_));
 sky130_fd_sc_hd__a22o_1 _6596_ (.A1(net368),
    .A2(net315),
    .B1(net257),
    .B2(net892),
    .X(_0921_));
 sky130_fd_sc_hd__or2_4 _6597_ (.A(_1283_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .X(_3416_));
 sky130_fd_sc_hd__nor3_2 _6598_ (.A(_2613_),
    .B(_2614_),
    .C(_3416_),
    .Y(_3417_));
 sky130_fd_sc_hd__or3_4 _6599_ (.A(_2613_),
    .B(_2614_),
    .C(_3416_),
    .X(_3418_));
 sky130_fd_sc_hd__and2_1 _6600_ (.A(net329),
    .B(net313),
    .X(_3419_));
 sky130_fd_sc_hd__a31o_1 _6601_ (.A1(net462),
    .A2(net1798),
    .A3(net311),
    .B1(_3419_),
    .X(_0922_));
 sky130_fd_sc_hd__and2_1 _6602_ (.A(net330),
    .B(net313),
    .X(_3420_));
 sky130_fd_sc_hd__a31o_1 _6603_ (.A1(net460),
    .A2(net1802),
    .A3(net311),
    .B1(_3420_),
    .X(_0923_));
 sky130_fd_sc_hd__or3_1 _6604_ (.A(net472),
    .B(net2093),
    .C(net313),
    .X(_3421_));
 sky130_fd_sc_hd__o21a_1 _6605_ (.A1(net331),
    .A2(net311),
    .B1(_3421_),
    .X(_0924_));
 sky130_fd_sc_hd__and2_1 _6606_ (.A(net332),
    .B(net313),
    .X(_3422_));
 sky130_fd_sc_hd__a31o_1 _6607_ (.A1(net462),
    .A2(net1824),
    .A3(_3418_),
    .B1(_3422_),
    .X(_0925_));
 sky130_fd_sc_hd__and2_1 _6608_ (.A(net327),
    .B(net313),
    .X(_3423_));
 sky130_fd_sc_hd__a31o_1 _6609_ (.A1(net459),
    .A2(net1800),
    .A3(net311),
    .B1(_3423_),
    .X(_0926_));
 sky130_fd_sc_hd__nor2_1 _6610_ (.A(_1607_),
    .B(net311),
    .Y(_3424_));
 sky130_fd_sc_hd__a31o_1 _6611_ (.A1(net458),
    .A2(net1893),
    .A3(net311),
    .B1(_3424_),
    .X(_0927_));
 sky130_fd_sc_hd__and2_1 _6612_ (.A(net326),
    .B(net313),
    .X(_3425_));
 sky130_fd_sc_hd__a31o_1 _6613_ (.A1(net456),
    .A2(net1840),
    .A3(net311),
    .B1(_3425_),
    .X(_0928_));
 sky130_fd_sc_hd__and2_1 _6614_ (.A(net328),
    .B(net313),
    .X(_3426_));
 sky130_fd_sc_hd__a31o_1 _6615_ (.A1(net455),
    .A2(net1830),
    .A3(net311),
    .B1(_3426_),
    .X(_0929_));
 sky130_fd_sc_hd__and2_1 _6616_ (.A(net323),
    .B(net312),
    .X(_3427_));
 sky130_fd_sc_hd__a31o_1 _6617_ (.A1(net458),
    .A2(net1916),
    .A3(net311),
    .B1(_3427_),
    .X(_0930_));
 sky130_fd_sc_hd__and2_1 _6618_ (.A(net325),
    .B(net313),
    .X(_3428_));
 sky130_fd_sc_hd__a31o_1 _6619_ (.A1(net461),
    .A2(net1937),
    .A3(net311),
    .B1(_3428_),
    .X(_0931_));
 sky130_fd_sc_hd__and2_1 _6620_ (.A(net324),
    .B(net313),
    .X(_3429_));
 sky130_fd_sc_hd__a31o_1 _6621_ (.A1(net455),
    .A2(net1941),
    .A3(net311),
    .B1(_3429_),
    .X(_0932_));
 sky130_fd_sc_hd__and2_1 _6622_ (.A(net322),
    .B(net312),
    .X(_3430_));
 sky130_fd_sc_hd__a31o_1 _6623_ (.A1(net447),
    .A2(net1876),
    .A3(net310),
    .B1(_3430_),
    .X(_0933_));
 sky130_fd_sc_hd__and2_1 _6624_ (.A(net319),
    .B(net313),
    .X(_3431_));
 sky130_fd_sc_hd__a31o_1 _6625_ (.A1(net459),
    .A2(net1950),
    .A3(net311),
    .B1(_3431_),
    .X(_0934_));
 sky130_fd_sc_hd__and2_1 _6626_ (.A(net321),
    .B(net312),
    .X(_3432_));
 sky130_fd_sc_hd__a31o_1 _6627_ (.A1(net454),
    .A2(net1746),
    .A3(net310),
    .B1(_3432_),
    .X(_0935_));
 sky130_fd_sc_hd__and2_1 _6628_ (.A(net320),
    .B(net312),
    .X(_3433_));
 sky130_fd_sc_hd__a31o_1 _6629_ (.A1(net452),
    .A2(net1838),
    .A3(_3418_),
    .B1(_3433_),
    .X(_0936_));
 sky130_fd_sc_hd__and2_1 _6630_ (.A(net318),
    .B(net313),
    .X(_3434_));
 sky130_fd_sc_hd__a31o_1 _6631_ (.A1(net458),
    .A2(net1812),
    .A3(net311),
    .B1(_3434_),
    .X(_0937_));
 sky130_fd_sc_hd__and2_1 _6632_ (.A(net342),
    .B(net312),
    .X(_3435_));
 sky130_fd_sc_hd__a31o_1 _6633_ (.A1(net454),
    .A2(net1891),
    .A3(net310),
    .B1(_3435_),
    .X(_0938_));
 sky130_fd_sc_hd__nor2_1 _6634_ (.A(_1381_),
    .B(net310),
    .Y(_3436_));
 sky130_fd_sc_hd__a31o_1 _6635_ (.A1(net445),
    .A2(net1866),
    .A3(net310),
    .B1(_3436_),
    .X(_0939_));
 sky130_fd_sc_hd__and2_1 _6636_ (.A(net341),
    .B(net313),
    .X(_3437_));
 sky130_fd_sc_hd__a31o_1 _6637_ (.A1(net460),
    .A2(net1851),
    .A3(net311),
    .B1(_3437_),
    .X(_0940_));
 sky130_fd_sc_hd__and2_1 _6638_ (.A(net343),
    .B(net312),
    .X(_3438_));
 sky130_fd_sc_hd__a31o_1 _6639_ (.A1(net450),
    .A2(net1730),
    .A3(net310),
    .B1(_3438_),
    .X(_0941_));
 sky130_fd_sc_hd__and2_1 _6640_ (.A(net338),
    .B(net312),
    .X(_3439_));
 sky130_fd_sc_hd__a31o_1 _6641_ (.A1(net445),
    .A2(net1834),
    .A3(net310),
    .B1(_3439_),
    .X(_0942_));
 sky130_fd_sc_hd__and2_1 _6642_ (.A(net340),
    .B(net312),
    .X(_3440_));
 sky130_fd_sc_hd__a31o_1 _6643_ (.A1(net445),
    .A2(net1846),
    .A3(net310),
    .B1(_3440_),
    .X(_0943_));
 sky130_fd_sc_hd__and2_1 _6644_ (.A(net339),
    .B(net312),
    .X(_3441_));
 sky130_fd_sc_hd__a31o_1 _6645_ (.A1(net453),
    .A2(net1963),
    .A3(net310),
    .B1(_3441_),
    .X(_0944_));
 sky130_fd_sc_hd__and2_1 _6646_ (.A(net337),
    .B(net312),
    .X(_3442_));
 sky130_fd_sc_hd__a31o_1 _6647_ (.A1(net446),
    .A2(net1895),
    .A3(net310),
    .B1(_3442_),
    .X(_0945_));
 sky130_fd_sc_hd__and2_1 _6648_ (.A(net334),
    .B(net313),
    .X(_3443_));
 sky130_fd_sc_hd__a31o_1 _6649_ (.A1(net461),
    .A2(net1781),
    .A3(net311),
    .B1(_3443_),
    .X(_0946_));
 sky130_fd_sc_hd__and2_1 _6650_ (.A(net336),
    .B(net312),
    .X(_3444_));
 sky130_fd_sc_hd__a31o_1 _6651_ (.A1(net446),
    .A2(net1910),
    .A3(net310),
    .B1(_3444_),
    .X(_0947_));
 sky130_fd_sc_hd__and2_1 _6652_ (.A(net335),
    .B(net312),
    .X(_3445_));
 sky130_fd_sc_hd__a31o_1 _6653_ (.A1(net446),
    .A2(net1929),
    .A3(net310),
    .B1(_3445_),
    .X(_0948_));
 sky130_fd_sc_hd__and2_1 _6654_ (.A(net333),
    .B(net312),
    .X(_3446_));
 sky130_fd_sc_hd__a31o_1 _6655_ (.A1(net454),
    .A2(net1908),
    .A3(net310),
    .B1(_3446_),
    .X(_0949_));
 sky130_fd_sc_hd__and2_1 _6656_ (.A(net346),
    .B(net312),
    .X(_3447_));
 sky130_fd_sc_hd__a31o_1 _6657_ (.A1(net447),
    .A2(net1897),
    .A3(net310),
    .B1(_3447_),
    .X(_0950_));
 sky130_fd_sc_hd__and2_1 _6658_ (.A(net344),
    .B(net312),
    .X(_3448_));
 sky130_fd_sc_hd__a31o_1 _6659_ (.A1(net445),
    .A2(net1785),
    .A3(net310),
    .B1(_3448_),
    .X(_0951_));
 sky130_fd_sc_hd__and2_1 _6660_ (.A(net345),
    .B(net313),
    .X(_3449_));
 sky130_fd_sc_hd__a31o_1 _6661_ (.A1(net461),
    .A2(net1906),
    .A3(net311),
    .B1(_3449_),
    .X(_0952_));
 sky130_fd_sc_hd__and2_1 _6662_ (.A(net368),
    .B(net312),
    .X(_3450_));
 sky130_fd_sc_hd__a31o_1 _6663_ (.A1(net448),
    .A2(net1768),
    .A3(net310),
    .B1(_3450_),
    .X(_0953_));
 sky130_fd_sc_hd__nor2_2 _6664_ (.A(_2628_),
    .B(_3416_),
    .Y(_3451_));
 sky130_fd_sc_hd__or2_1 _6665_ (.A(_2628_),
    .B(_3416_),
    .X(_3452_));
 sky130_fd_sc_hd__nor2_2 _6666_ (.A(net471),
    .B(net256),
    .Y(_3453_));
 sky130_fd_sc_hd__nand2_1 _6667_ (.A(net462),
    .B(_3452_),
    .Y(_3454_));
 sky130_fd_sc_hd__o22a_1 _6668_ (.A1(net329),
    .A2(_3452_),
    .B1(_3454_),
    .B2(net805),
    .X(_0954_));
 sky130_fd_sc_hd__a22o_1 _6669_ (.A1(net330),
    .A2(net256),
    .B1(net220),
    .B2(net1456),
    .X(_0955_));
 sky130_fd_sc_hd__o22a_1 _6670_ (.A1(net331),
    .A2(_3452_),
    .B1(_3454_),
    .B2(net794),
    .X(_0956_));
 sky130_fd_sc_hd__a22o_1 _6671_ (.A1(net332),
    .A2(net256),
    .B1(net220),
    .B2(net1071),
    .X(_0957_));
 sky130_fd_sc_hd__a22o_1 _6672_ (.A1(net327),
    .A2(net256),
    .B1(net220),
    .B2(net1504),
    .X(_0958_));
 sky130_fd_sc_hd__a22o_1 _6673_ (.A1(_1608_),
    .A2(net256),
    .B1(net220),
    .B2(net1075),
    .X(_0959_));
 sky130_fd_sc_hd__a22o_1 _6674_ (.A1(net326),
    .A2(net256),
    .B1(net220),
    .B2(net1203),
    .X(_0960_));
 sky130_fd_sc_hd__a22o_1 _6675_ (.A1(net328),
    .A2(net256),
    .B1(net220),
    .B2(net1444),
    .X(_0961_));
 sky130_fd_sc_hd__a22o_1 _6676_ (.A1(net323),
    .A2(net256),
    .B1(net220),
    .B2(net1187),
    .X(_0962_));
 sky130_fd_sc_hd__a22o_1 _6677_ (.A1(net325),
    .A2(net256),
    .B1(net220),
    .B2(net1173),
    .X(_0963_));
 sky130_fd_sc_hd__a22o_1 _6678_ (.A1(net324),
    .A2(net256),
    .B1(net220),
    .B2(net1678),
    .X(_0964_));
 sky130_fd_sc_hd__a22o_1 _6679_ (.A1(net322),
    .A2(net255),
    .B1(net219),
    .B2(net1019),
    .X(_0965_));
 sky130_fd_sc_hd__a22o_1 _6680_ (.A1(net319),
    .A2(net256),
    .B1(net220),
    .B2(net1586),
    .X(_0966_));
 sky130_fd_sc_hd__a22o_1 _6681_ (.A1(net321),
    .A2(net255),
    .B1(net219),
    .B2(net1127),
    .X(_0967_));
 sky130_fd_sc_hd__a22o_1 _6682_ (.A1(net320),
    .A2(net255),
    .B1(net219),
    .B2(net1371),
    .X(_0968_));
 sky130_fd_sc_hd__a22o_1 _6683_ (.A1(net318),
    .A2(net256),
    .B1(net220),
    .B2(net1035),
    .X(_0969_));
 sky130_fd_sc_hd__a22o_1 _6684_ (.A1(net342),
    .A2(net255),
    .B1(net219),
    .B2(net1498),
    .X(_0970_));
 sky130_fd_sc_hd__a22o_1 _6685_ (.A1(_1382_),
    .A2(net255),
    .B1(net219),
    .B2(net1221),
    .X(_0971_));
 sky130_fd_sc_hd__a22o_1 _6686_ (.A1(net341),
    .A2(net256),
    .B1(net220),
    .B2(net1484),
    .X(_0972_));
 sky130_fd_sc_hd__a22o_1 _6687_ (.A1(net343),
    .A2(net255),
    .B1(net219),
    .B2(net1007),
    .X(_0973_));
 sky130_fd_sc_hd__a22o_1 _6688_ (.A1(net338),
    .A2(net255),
    .B1(net219),
    .B2(net1207),
    .X(_0974_));
 sky130_fd_sc_hd__a22o_1 _6689_ (.A1(net340),
    .A2(net255),
    .B1(net219),
    .B2(net1566),
    .X(_0975_));
 sky130_fd_sc_hd__a22o_1 _6690_ (.A1(net339),
    .A2(net255),
    .B1(net219),
    .B2(net1588),
    .X(_0976_));
 sky130_fd_sc_hd__a22o_1 _6691_ (.A1(net337),
    .A2(net255),
    .B1(net219),
    .B2(net1309),
    .X(_0977_));
 sky130_fd_sc_hd__a22o_1 _6692_ (.A1(net334),
    .A2(net256),
    .B1(net220),
    .B2(net979),
    .X(_0978_));
 sky130_fd_sc_hd__a22o_1 _6693_ (.A1(net336),
    .A2(net255),
    .B1(net219),
    .B2(net1568),
    .X(_0979_));
 sky130_fd_sc_hd__a22o_1 _6694_ (.A1(net335),
    .A2(net255),
    .B1(net219),
    .B2(net1752),
    .X(_0980_));
 sky130_fd_sc_hd__a22o_1 _6695_ (.A1(net333),
    .A2(net255),
    .B1(net219),
    .B2(net1454),
    .X(_0981_));
 sky130_fd_sc_hd__a22o_1 _6696_ (.A1(net346),
    .A2(net255),
    .B1(net219),
    .B2(net981),
    .X(_0982_));
 sky130_fd_sc_hd__a22o_1 _6697_ (.A1(net344),
    .A2(net255),
    .B1(net219),
    .B2(net1490),
    .X(_0983_));
 sky130_fd_sc_hd__a22o_1 _6698_ (.A1(net345),
    .A2(net256),
    .B1(net220),
    .B2(net1121),
    .X(_0984_));
 sky130_fd_sc_hd__a22o_1 _6699_ (.A1(net368),
    .A2(net255),
    .B1(net219),
    .B2(net1701),
    .X(_0985_));
 sky130_fd_sc_hd__or2_2 _6700_ (.A(_2614_),
    .B(_2623_),
    .X(_3455_));
 sky130_fd_sc_hd__nor2_2 _6701_ (.A(_2637_),
    .B(_3455_),
    .Y(_3456_));
 sky130_fd_sc_hd__or2_2 _6702_ (.A(_2637_),
    .B(_3455_),
    .X(_3457_));
 sky130_fd_sc_hd__nor2_2 _6703_ (.A(net471),
    .B(net254),
    .Y(_3458_));
 sky130_fd_sc_hd__nand2_1 _6704_ (.A(net460),
    .B(_3457_),
    .Y(_3459_));
 sky130_fd_sc_hd__o22a_1 _6705_ (.A1(net329),
    .A2(_3457_),
    .B1(_3459_),
    .B2(net911),
    .X(_0986_));
 sky130_fd_sc_hd__o22a_1 _6706_ (.A1(net330),
    .A2(_3457_),
    .B1(_3459_),
    .B2(net1295),
    .X(_0987_));
 sky130_fd_sc_hd__a22o_1 _6707_ (.A1(net331),
    .A2(net254),
    .B1(net218),
    .B2(net1199),
    .X(_0988_));
 sky130_fd_sc_hd__o22a_1 _6708_ (.A1(net332),
    .A2(_3457_),
    .B1(_3459_),
    .B2(net867),
    .X(_0989_));
 sky130_fd_sc_hd__a22o_1 _6709_ (.A1(net327),
    .A2(net254),
    .B1(net218),
    .B2(net1436),
    .X(_0990_));
 sky130_fd_sc_hd__a22o_1 _6710_ (.A1(_1608_),
    .A2(net254),
    .B1(net218),
    .B2(net1335),
    .X(_0991_));
 sky130_fd_sc_hd__a22o_1 _6711_ (.A1(net326),
    .A2(net254),
    .B1(net218),
    .B2(net1009),
    .X(_0992_));
 sky130_fd_sc_hd__a22o_1 _6712_ (.A1(net328),
    .A2(net253),
    .B1(net217),
    .B2(net1405),
    .X(_0993_));
 sky130_fd_sc_hd__a22o_1 _6713_ (.A1(net323),
    .A2(net254),
    .B1(net218),
    .B2(net1205),
    .X(_0994_));
 sky130_fd_sc_hd__a22o_1 _6714_ (.A1(net325),
    .A2(net254),
    .B1(net218),
    .B2(net1237),
    .X(_0995_));
 sky130_fd_sc_hd__a22o_1 _6715_ (.A1(net324),
    .A2(net254),
    .B1(net218),
    .B2(net1383),
    .X(_0996_));
 sky130_fd_sc_hd__a22o_1 _6716_ (.A1(net322),
    .A2(net253),
    .B1(net217),
    .B2(net1185),
    .X(_0997_));
 sky130_fd_sc_hd__a22o_1 _6717_ (.A1(net319),
    .A2(net254),
    .B1(net218),
    .B2(net1393),
    .X(_0998_));
 sky130_fd_sc_hd__a22o_1 _6718_ (.A1(net321),
    .A2(net253),
    .B1(net217),
    .B2(net1592),
    .X(_0999_));
 sky130_fd_sc_hd__a22o_1 _6719_ (.A1(net320),
    .A2(net253),
    .B1(net217),
    .B2(net1576),
    .X(_1000_));
 sky130_fd_sc_hd__a22o_1 _6720_ (.A1(net318),
    .A2(net254),
    .B1(net218),
    .B2(net1385),
    .X(_1001_));
 sky130_fd_sc_hd__a22o_1 _6721_ (.A1(net342),
    .A2(net253),
    .B1(net217),
    .B2(net1438),
    .X(_1002_));
 sky130_fd_sc_hd__a22o_1 _6722_ (.A1(_1382_),
    .A2(net253),
    .B1(net217),
    .B2(net1415),
    .X(_1003_));
 sky130_fd_sc_hd__a22o_1 _6723_ (.A1(net341),
    .A2(net254),
    .B1(net218),
    .B2(net1277),
    .X(_1004_));
 sky130_fd_sc_hd__a22o_1 _6724_ (.A1(net343),
    .A2(net253),
    .B1(net217),
    .B2(net927),
    .X(_1005_));
 sky130_fd_sc_hd__a22o_1 _6725_ (.A1(net338),
    .A2(net253),
    .B1(net217),
    .B2(net1540),
    .X(_1006_));
 sky130_fd_sc_hd__a22o_1 _6726_ (.A1(net340),
    .A2(net253),
    .B1(net217),
    .B2(net1756),
    .X(_1007_));
 sky130_fd_sc_hd__a22o_1 _6727_ (.A1(net339),
    .A2(net254),
    .B1(net218),
    .B2(net1273),
    .X(_1008_));
 sky130_fd_sc_hd__a22o_1 _6728_ (.A1(net337),
    .A2(net253),
    .B1(net217),
    .B2(net1460),
    .X(_1009_));
 sky130_fd_sc_hd__a22o_1 _6729_ (.A1(net334),
    .A2(net254),
    .B1(net218),
    .B2(net1343),
    .X(_1010_));
 sky130_fd_sc_hd__a22o_1 _6730_ (.A1(net336),
    .A2(net253),
    .B1(net217),
    .B2(net1397),
    .X(_1011_));
 sky130_fd_sc_hd__a22o_1 _6731_ (.A1(net335),
    .A2(net253),
    .B1(net217),
    .B2(net1560),
    .X(_1012_));
 sky130_fd_sc_hd__a22o_1 _6732_ (.A1(net333),
    .A2(net253),
    .B1(net217),
    .B2(net1045),
    .X(_1013_));
 sky130_fd_sc_hd__a22o_1 _6733_ (.A1(net346),
    .A2(net253),
    .B1(net217),
    .B2(net1161),
    .X(_1014_));
 sky130_fd_sc_hd__a22o_1 _6734_ (.A1(net344),
    .A2(net253),
    .B1(net217),
    .B2(net1211),
    .X(_1015_));
 sky130_fd_sc_hd__a22o_1 _6735_ (.A1(net345),
    .A2(net254),
    .B1(net218),
    .B2(net1005),
    .X(_1016_));
 sky130_fd_sc_hd__a22o_1 _6736_ (.A1(net368),
    .A2(net253),
    .B1(net217),
    .B2(net1191),
    .X(_1017_));
 sky130_fd_sc_hd__nor2_2 _6737_ (.A(_2613_),
    .B(_3455_),
    .Y(_3460_));
 sky130_fd_sc_hd__or2_4 _6738_ (.A(_2613_),
    .B(_3455_),
    .X(_3461_));
 sky130_fd_sc_hd__and2_1 _6739_ (.A(net329),
    .B(net252),
    .X(_3462_));
 sky130_fd_sc_hd__a31o_1 _6740_ (.A1(net460),
    .A2(net1931),
    .A3(net249),
    .B1(_3462_),
    .X(_1018_));
 sky130_fd_sc_hd__and2_1 _6741_ (.A(net330),
    .B(net252),
    .X(_3463_));
 sky130_fd_sc_hd__a31o_1 _6742_ (.A1(net462),
    .A2(net1818),
    .A3(net249),
    .B1(_3463_),
    .X(_1019_));
 sky130_fd_sc_hd__and2_1 _6743_ (.A(net331),
    .B(net252),
    .X(_3464_));
 sky130_fd_sc_hd__a31o_1 _6744_ (.A1(net456),
    .A2(net1684),
    .A3(net249),
    .B1(_3464_),
    .X(_1020_));
 sky130_fd_sc_hd__or3_1 _6745_ (.A(net471),
    .B(net2102),
    .C(net251),
    .X(_3465_));
 sky130_fd_sc_hd__o21a_1 _6746_ (.A1(_1523_),
    .A2(net249),
    .B1(_3465_),
    .X(_1021_));
 sky130_fd_sc_hd__and2_1 _6747_ (.A(net327),
    .B(net252),
    .X(_3466_));
 sky130_fd_sc_hd__a31o_1 _6748_ (.A1(net459),
    .A2(net1980),
    .A3(net249),
    .B1(_3466_),
    .X(_1022_));
 sky130_fd_sc_hd__nor2_1 _6749_ (.A(_1607_),
    .B(net249),
    .Y(_3467_));
 sky130_fd_sc_hd__a31o_1 _6750_ (.A1(net458),
    .A2(net1762),
    .A3(net249),
    .B1(_3467_),
    .X(_1023_));
 sky130_fd_sc_hd__and2_1 _6751_ (.A(net326),
    .B(net252),
    .X(_3468_));
 sky130_fd_sc_hd__a31o_1 _6752_ (.A1(net456),
    .A2(net1870),
    .A3(net249),
    .B1(_3468_),
    .X(_1024_));
 sky130_fd_sc_hd__and2_1 _6753_ (.A(net328),
    .B(net251),
    .X(_3469_));
 sky130_fd_sc_hd__a31o_1 _6754_ (.A1(net455),
    .A2(net1899),
    .A3(net250),
    .B1(_3469_),
    .X(_1025_));
 sky130_fd_sc_hd__and2_1 _6755_ (.A(net323),
    .B(net252),
    .X(_3470_));
 sky130_fd_sc_hd__a31o_1 _6756_ (.A1(net452),
    .A2(net1948),
    .A3(net249),
    .B1(_3470_),
    .X(_1026_));
 sky130_fd_sc_hd__and2_1 _6757_ (.A(net325),
    .B(net252),
    .X(_3471_));
 sky130_fd_sc_hd__a31o_1 _6758_ (.A1(net461),
    .A2(net1709),
    .A3(_3461_),
    .B1(_3471_),
    .X(_1027_));
 sky130_fd_sc_hd__and2_1 _6759_ (.A(net324),
    .B(net252),
    .X(_3472_));
 sky130_fd_sc_hd__a31o_1 _6760_ (.A1(net460),
    .A2(net1772),
    .A3(_3461_),
    .B1(_3472_),
    .X(_1028_));
 sky130_fd_sc_hd__and2_1 _6761_ (.A(net322),
    .B(net251),
    .X(_3473_));
 sky130_fd_sc_hd__a31o_1 _6762_ (.A1(net447),
    .A2(net1858),
    .A3(net250),
    .B1(_3473_),
    .X(_1029_));
 sky130_fd_sc_hd__and2_1 _6763_ (.A(net319),
    .B(net252),
    .X(_3474_));
 sky130_fd_sc_hd__a31o_1 _6764_ (.A1(net459),
    .A2(net1926),
    .A3(net249),
    .B1(_3474_),
    .X(_1030_));
 sky130_fd_sc_hd__and2_1 _6765_ (.A(net321),
    .B(net251),
    .X(_3475_));
 sky130_fd_sc_hd__a31o_1 _6766_ (.A1(net454),
    .A2(net1860),
    .A3(net250),
    .B1(_3475_),
    .X(_1031_));
 sky130_fd_sc_hd__and2_1 _6767_ (.A(net320),
    .B(net251),
    .X(_3476_));
 sky130_fd_sc_hd__a31o_1 _6768_ (.A1(net452),
    .A2(net1956),
    .A3(net249),
    .B1(_3476_),
    .X(_1032_));
 sky130_fd_sc_hd__and2_1 _6769_ (.A(net318),
    .B(net252),
    .X(_3477_));
 sky130_fd_sc_hd__a31o_1 _6770_ (.A1(net458),
    .A2(net1622),
    .A3(net249),
    .B1(_3477_),
    .X(_1033_));
 sky130_fd_sc_hd__and2_1 _6771_ (.A(net342),
    .B(net251),
    .X(_3478_));
 sky130_fd_sc_hd__a31o_1 _6772_ (.A1(net453),
    .A2(net1662),
    .A3(net250),
    .B1(_3478_),
    .X(_1034_));
 sky130_fd_sc_hd__nor2_1 _6773_ (.A(_1381_),
    .B(net250),
    .Y(_3479_));
 sky130_fd_sc_hd__a31o_1 _6774_ (.A1(net447),
    .A2(net1902),
    .A3(net250),
    .B1(_3479_),
    .X(_1035_));
 sky130_fd_sc_hd__and2_1 _6775_ (.A(net341),
    .B(net252),
    .X(_3480_));
 sky130_fd_sc_hd__a31o_1 _6776_ (.A1(net460),
    .A2(net1820),
    .A3(net249),
    .B1(_3480_),
    .X(_1036_));
 sky130_fd_sc_hd__and2_1 _6777_ (.A(net343),
    .B(net251),
    .X(_3481_));
 sky130_fd_sc_hd__a31o_1 _6778_ (.A1(net450),
    .A2(net1734),
    .A3(net250),
    .B1(_3481_),
    .X(_1037_));
 sky130_fd_sc_hd__and2_1 _6779_ (.A(_1452_),
    .B(net251),
    .X(_3482_));
 sky130_fd_sc_hd__a31o_1 _6780_ (.A1(net445),
    .A2(net1883),
    .A3(net250),
    .B1(_3482_),
    .X(_1038_));
 sky130_fd_sc_hd__and2_1 _6781_ (.A(net340),
    .B(net251),
    .X(_3483_));
 sky130_fd_sc_hd__a31o_1 _6782_ (.A1(net448),
    .A2(net1776),
    .A3(net250),
    .B1(_3483_),
    .X(_1039_));
 sky130_fd_sc_hd__and2_1 _6783_ (.A(net339),
    .B(net252),
    .X(_3484_));
 sky130_fd_sc_hd__a31o_1 _6784_ (.A1(net455),
    .A2(net1965),
    .A3(net249),
    .B1(_3484_),
    .X(_1040_));
 sky130_fd_sc_hd__and2_1 _6785_ (.A(net337),
    .B(net251),
    .X(_3485_));
 sky130_fd_sc_hd__a31o_1 _6786_ (.A1(net446),
    .A2(net1922),
    .A3(net250),
    .B1(_3485_),
    .X(_1041_));
 sky130_fd_sc_hd__and2_1 _6787_ (.A(net334),
    .B(net252),
    .X(_3486_));
 sky130_fd_sc_hd__a31o_1 _6788_ (.A1(net461),
    .A2(net1924),
    .A3(net249),
    .B1(_3486_),
    .X(_1042_));
 sky130_fd_sc_hd__and2_1 _6789_ (.A(net336),
    .B(net251),
    .X(_3487_));
 sky130_fd_sc_hd__a31o_1 _6790_ (.A1(net446),
    .A2(net1914),
    .A3(net250),
    .B1(_3487_),
    .X(_1043_));
 sky130_fd_sc_hd__and2_1 _6791_ (.A(net335),
    .B(net251),
    .X(_3488_));
 sky130_fd_sc_hd__a31o_1 _6792_ (.A1(net445),
    .A2(net1912),
    .A3(net250),
    .B1(_3488_),
    .X(_1044_));
 sky130_fd_sc_hd__and2_1 _6793_ (.A(net333),
    .B(net251),
    .X(_3489_));
 sky130_fd_sc_hd__a31o_1 _6794_ (.A1(net456),
    .A2(net1764),
    .A3(net250),
    .B1(_3489_),
    .X(_1045_));
 sky130_fd_sc_hd__and2_1 _6795_ (.A(net346),
    .B(net251),
    .X(_3490_));
 sky130_fd_sc_hd__a31o_1 _6796_ (.A1(net447),
    .A2(net1889),
    .A3(net250),
    .B1(_3490_),
    .X(_1046_));
 sky130_fd_sc_hd__and2_1 _6797_ (.A(net344),
    .B(net251),
    .X(_3491_));
 sky130_fd_sc_hd__a31o_1 _6798_ (.A1(net445),
    .A2(net1978),
    .A3(net250),
    .B1(_3491_),
    .X(_1047_));
 sky130_fd_sc_hd__and2_1 _6799_ (.A(net345),
    .B(net252),
    .X(_3492_));
 sky130_fd_sc_hd__a31o_1 _6800_ (.A1(net461),
    .A2(net1795),
    .A3(net249),
    .B1(_3492_),
    .X(_1048_));
 sky130_fd_sc_hd__and2_1 _6801_ (.A(net368),
    .B(net251),
    .X(_3493_));
 sky130_fd_sc_hd__a31o_1 _6802_ (.A1(net447),
    .A2(net1705),
    .A3(net250),
    .B1(_3493_),
    .X(_1049_));
 sky130_fd_sc_hd__nor3_4 _6803_ (.A(_2614_),
    .B(_2637_),
    .C(_3416_),
    .Y(_3494_));
 sky130_fd_sc_hd__or3_2 _6804_ (.A(_2614_),
    .B(_2637_),
    .C(_3416_),
    .X(_3495_));
 sky130_fd_sc_hd__nor2_4 _6805_ (.A(net471),
    .B(net309),
    .Y(_3496_));
 sky130_fd_sc_hd__nand2_1 _6806_ (.A(net462),
    .B(_3495_),
    .Y(_3497_));
 sky130_fd_sc_hd__o22a_1 _6807_ (.A1(net329),
    .A2(_3495_),
    .B1(_3497_),
    .B2(net784),
    .X(_1050_));
 sky130_fd_sc_hd__o22a_1 _6808_ (.A1(net330),
    .A2(_3495_),
    .B1(_3497_),
    .B2(net1808),
    .X(_1051_));
 sky130_fd_sc_hd__o22a_1 _6809_ (.A1(net331),
    .A2(_3495_),
    .B1(_3497_),
    .B2(net797),
    .X(_1052_));
 sky130_fd_sc_hd__a22o_1 _6810_ (.A1(net332),
    .A2(net309),
    .B1(net248),
    .B2(net1470),
    .X(_1053_));
 sky130_fd_sc_hd__a22o_1 _6811_ (.A1(net327),
    .A2(net309),
    .B1(net248),
    .B2(net1387),
    .X(_1054_));
 sky130_fd_sc_hd__a22o_1 _6812_ (.A1(_1608_),
    .A2(net309),
    .B1(net248),
    .B2(net1089),
    .X(_1055_));
 sky130_fd_sc_hd__a22o_1 _6813_ (.A1(net326),
    .A2(net309),
    .B1(net248),
    .B2(net1259),
    .X(_1056_));
 sky130_fd_sc_hd__a22o_1 _6814_ (.A1(net328),
    .A2(net309),
    .B1(net248),
    .B2(net1532),
    .X(_1057_));
 sky130_fd_sc_hd__a22o_1 _6815_ (.A1(net323),
    .A2(net309),
    .B1(net248),
    .B2(net1428),
    .X(_1058_));
 sky130_fd_sc_hd__a22o_1 _6816_ (.A1(net325),
    .A2(net309),
    .B1(net248),
    .B2(net1157),
    .X(_1059_));
 sky130_fd_sc_hd__a22o_1 _6817_ (.A1(net324),
    .A2(net309),
    .B1(net248),
    .B2(net1452),
    .X(_1060_));
 sky130_fd_sc_hd__a22o_1 _6818_ (.A1(net322),
    .A2(net308),
    .B1(net247),
    .B2(net1508),
    .X(_1061_));
 sky130_fd_sc_hd__a22o_1 _6819_ (.A1(net319),
    .A2(net309),
    .B1(net248),
    .B2(net1548),
    .X(_1062_));
 sky130_fd_sc_hd__a22o_1 _6820_ (.A1(net321),
    .A2(net308),
    .B1(net247),
    .B2(net1375),
    .X(_1063_));
 sky130_fd_sc_hd__a22o_1 _6821_ (.A1(net320),
    .A2(net308),
    .B1(net247),
    .B2(net1079),
    .X(_1064_));
 sky130_fd_sc_hd__a22o_1 _6822_ (.A1(net318),
    .A2(net309),
    .B1(net248),
    .B2(net1241),
    .X(_1065_));
 sky130_fd_sc_hd__a22o_1 _6823_ (.A1(net342),
    .A2(net308),
    .B1(net247),
    .B2(net963),
    .X(_1066_));
 sky130_fd_sc_hd__a22o_1 _6824_ (.A1(_1382_),
    .A2(net308),
    .B1(net247),
    .B2(net907),
    .X(_1067_));
 sky130_fd_sc_hd__a22o_1 _6825_ (.A1(net341),
    .A2(net309),
    .B1(net248),
    .B2(net1492),
    .X(_1068_));
 sky130_fd_sc_hd__a22o_1 _6826_ (.A1(net343),
    .A2(net308),
    .B1(net247),
    .B2(net993),
    .X(_1069_));
 sky130_fd_sc_hd__a22o_1 _6827_ (.A1(net338),
    .A2(net308),
    .B1(net247),
    .B2(net1422),
    .X(_1070_));
 sky130_fd_sc_hd__a22o_1 _6828_ (.A1(net340),
    .A2(net308),
    .B1(net247),
    .B2(net1333),
    .X(_1071_));
 sky130_fd_sc_hd__a22o_1 _6829_ (.A1(net339),
    .A2(net308),
    .B1(net247),
    .B2(net1626),
    .X(_1072_));
 sky130_fd_sc_hd__a22o_1 _6830_ (.A1(net337),
    .A2(net308),
    .B1(net247),
    .B2(net1574),
    .X(_1073_));
 sky130_fd_sc_hd__a22o_1 _6831_ (.A1(net334),
    .A2(net309),
    .B1(net248),
    .B2(net973),
    .X(_1074_));
 sky130_fd_sc_hd__a22o_1 _6832_ (.A1(net336),
    .A2(net308),
    .B1(net247),
    .B2(net1688),
    .X(_1075_));
 sky130_fd_sc_hd__a22o_1 _6833_ (.A1(net335),
    .A2(net308),
    .B1(net247),
    .B2(net1536),
    .X(_1076_));
 sky130_fd_sc_hd__a22o_1 _6834_ (.A1(net333),
    .A2(net308),
    .B1(net247),
    .B2(net1434),
    .X(_1077_));
 sky130_fd_sc_hd__a22o_1 _6835_ (.A1(net346),
    .A2(net308),
    .B1(net247),
    .B2(net942),
    .X(_1078_));
 sky130_fd_sc_hd__a22o_1 _6836_ (.A1(net344),
    .A2(net308),
    .B1(net247),
    .B2(net1269),
    .X(_1079_));
 sky130_fd_sc_hd__a22o_1 _6837_ (.A1(net345),
    .A2(net309),
    .B1(net248),
    .B2(net1514),
    .X(_1080_));
 sky130_fd_sc_hd__a22o_1 _6838_ (.A1(net368),
    .A2(net308),
    .B1(net247),
    .B2(net985),
    .X(_1081_));
 sky130_fd_sc_hd__nor2_2 _6839_ (.A(_2622_),
    .B(_3416_),
    .Y(_3498_));
 sky130_fd_sc_hd__or2_1 _6840_ (.A(_2622_),
    .B(_3416_),
    .X(_3499_));
 sky130_fd_sc_hd__nor2_4 _6841_ (.A(net471),
    .B(net246),
    .Y(_3500_));
 sky130_fd_sc_hd__nand2_1 _6842_ (.A(net460),
    .B(_3499_),
    .Y(_3501_));
 sky130_fd_sc_hd__a22o_1 _6843_ (.A1(net329),
    .A2(net246),
    .B1(net216),
    .B2(net940),
    .X(_1082_));
 sky130_fd_sc_hd__o22a_1 _6844_ (.A1(net330),
    .A2(_3499_),
    .B1(_3501_),
    .B2(net1967),
    .X(_1083_));
 sky130_fd_sc_hd__o22a_1 _6845_ (.A1(net331),
    .A2(_3499_),
    .B1(_3501_),
    .B2(net786),
    .X(_1084_));
 sky130_fd_sc_hd__a22o_1 _6846_ (.A1(net332),
    .A2(net246),
    .B1(net216),
    .B2(net1315),
    .X(_1085_));
 sky130_fd_sc_hd__a22o_1 _6847_ (.A1(net327),
    .A2(net246),
    .B1(net216),
    .B2(net1305),
    .X(_1086_));
 sky130_fd_sc_hd__a22o_1 _6848_ (.A1(_1608_),
    .A2(net246),
    .B1(net216),
    .B2(net1389),
    .X(_1087_));
 sky130_fd_sc_hd__a22o_1 _6849_ (.A1(net326),
    .A2(net246),
    .B1(net216),
    .B2(net1363),
    .X(_1088_));
 sky130_fd_sc_hd__a22o_1 _6850_ (.A1(net328),
    .A2(net246),
    .B1(net215),
    .B2(net1243),
    .X(_1089_));
 sky130_fd_sc_hd__a22o_1 _6851_ (.A1(net323),
    .A2(net245),
    .B1(net216),
    .B2(net1359),
    .X(_1090_));
 sky130_fd_sc_hd__a22o_1 _6852_ (.A1(net325),
    .A2(net246),
    .B1(net216),
    .B2(net1486),
    .X(_1091_));
 sky130_fd_sc_hd__a22o_1 _6853_ (.A1(net324),
    .A2(net246),
    .B1(net216),
    .B2(net1524),
    .X(_1092_));
 sky130_fd_sc_hd__a22o_1 _6854_ (.A1(net322),
    .A2(net245),
    .B1(net215),
    .B2(net1297),
    .X(_1093_));
 sky130_fd_sc_hd__a22o_1 _6855_ (.A1(net319),
    .A2(net246),
    .B1(net216),
    .B2(net1141),
    .X(_1094_));
 sky130_fd_sc_hd__a22o_1 _6856_ (.A1(net321),
    .A2(net245),
    .B1(net215),
    .B2(net1109),
    .X(_1095_));
 sky130_fd_sc_hd__a22o_1 _6857_ (.A1(net320),
    .A2(net246),
    .B1(net216),
    .B2(net1311),
    .X(_1096_));
 sky130_fd_sc_hd__a22o_1 _6858_ (.A1(net318),
    .A2(net246),
    .B1(net216),
    .B2(net1301),
    .X(_1097_));
 sky130_fd_sc_hd__a22o_1 _6859_ (.A1(net342),
    .A2(net245),
    .B1(net215),
    .B2(net1143),
    .X(_1098_));
 sky130_fd_sc_hd__a22o_1 _6860_ (.A1(_1382_),
    .A2(net245),
    .B1(net215),
    .B2(net1225),
    .X(_1099_));
 sky130_fd_sc_hd__a22o_1 _6861_ (.A1(net341),
    .A2(net246),
    .B1(net216),
    .B2(net1530),
    .X(_1100_));
 sky130_fd_sc_hd__a22o_1 _6862_ (.A1(net343),
    .A2(net245),
    .B1(net215),
    .B2(net1027),
    .X(_1101_));
 sky130_fd_sc_hd__a22o_1 _6863_ (.A1(net338),
    .A2(net245),
    .B1(net215),
    .B2(net1081),
    .X(_1102_));
 sky130_fd_sc_hd__a22o_1 _6864_ (.A1(net340),
    .A2(net245),
    .B1(net215),
    .B2(net1137),
    .X(_1103_));
 sky130_fd_sc_hd__a22o_1 _6865_ (.A1(net339),
    .A2(net245),
    .B1(net215),
    .B2(net1648),
    .X(_1104_));
 sky130_fd_sc_hd__a22o_1 _6866_ (.A1(_1463_),
    .A2(net245),
    .B1(net215),
    .B2(net1163),
    .X(_1105_));
 sky130_fd_sc_hd__a22o_1 _6867_ (.A1(net334),
    .A2(net246),
    .B1(net216),
    .B2(net917),
    .X(_1106_));
 sky130_fd_sc_hd__a22o_1 _6868_ (.A1(net336),
    .A2(net245),
    .B1(net215),
    .B2(net1271),
    .X(_1107_));
 sky130_fd_sc_hd__a22o_1 _6869_ (.A1(net335),
    .A2(net245),
    .B1(net215),
    .B2(net1091),
    .X(_1108_));
 sky130_fd_sc_hd__a22o_1 _6870_ (.A1(net333),
    .A2(net245),
    .B1(net215),
    .B2(net944),
    .X(_1109_));
 sky130_fd_sc_hd__a22o_1 _6871_ (.A1(net346),
    .A2(net245),
    .B1(net215),
    .B2(net991),
    .X(_1110_));
 sky130_fd_sc_hd__a22o_1 _6872_ (.A1(net344),
    .A2(net245),
    .B1(net215),
    .B2(net1401),
    .X(_1111_));
 sky130_fd_sc_hd__a22o_1 _6873_ (.A1(net345),
    .A2(net246),
    .B1(net216),
    .B2(net1331),
    .X(_1112_));
 sky130_fd_sc_hd__a22o_1 _6874_ (.A1(net368),
    .A2(net245),
    .B1(net215),
    .B2(net932),
    .X(_1113_));
 sky130_fd_sc_hd__nor3_1 _6875_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2622_),
    .Y(_3502_));
 sky130_fd_sc_hd__or3_4 _6876_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2622_),
    .X(_3503_));
 sky130_fd_sc_hd__and2_1 _6877_ (.A(net329),
    .B(net243),
    .X(_3504_));
 sky130_fd_sc_hd__a31o_1 _6878_ (.A1(net462),
    .A2(net1952),
    .A3(net241),
    .B1(_3504_),
    .X(_1144_));
 sky130_fd_sc_hd__or3_1 _6879_ (.A(net471),
    .B(net2086),
    .C(net243),
    .X(_3505_));
 sky130_fd_sc_hd__o21a_1 _6880_ (.A1(net330),
    .A2(net241),
    .B1(_3505_),
    .X(_1145_));
 sky130_fd_sc_hd__and2_1 _6881_ (.A(net331),
    .B(net243),
    .X(_3506_));
 sky130_fd_sc_hd__a31o_1 _6882_ (.A1(net456),
    .A2(net1740),
    .A3(net241),
    .B1(_3506_),
    .X(_1146_));
 sky130_fd_sc_hd__and2_1 _6883_ (.A(net332),
    .B(net244),
    .X(_3507_));
 sky130_fd_sc_hd__a31o_1 _6884_ (.A1(net462),
    .A2(net1628),
    .A3(_3503_),
    .B1(_3507_),
    .X(_1147_));
 sky130_fd_sc_hd__and2_1 _6885_ (.A(net327),
    .B(net243),
    .X(_3508_));
 sky130_fd_sc_hd__a31o_1 _6886_ (.A1(net459),
    .A2(net1636),
    .A3(net241),
    .B1(_3508_),
    .X(_1148_));
 sky130_fd_sc_hd__or3b_1 _6887_ (.A(net470),
    .B(net243),
    .C_N(net2127),
    .X(_3509_));
 sky130_fd_sc_hd__o21ai_1 _6888_ (.A1(_1607_),
    .A2(net241),
    .B1(_3509_),
    .Y(_1149_));
 sky130_fd_sc_hd__and2_1 _6889_ (.A(net326),
    .B(net243),
    .X(_3510_));
 sky130_fd_sc_hd__a31o_1 _6890_ (.A1(net456),
    .A2(net1744),
    .A3(net241),
    .B1(_3510_),
    .X(_1150_));
 sky130_fd_sc_hd__and2_1 _6891_ (.A(net328),
    .B(net243),
    .X(_3511_));
 sky130_fd_sc_hd__a31o_1 _6892_ (.A1(net455),
    .A2(net1770),
    .A3(net241),
    .B1(_3511_),
    .X(_1151_));
 sky130_fd_sc_hd__and2_1 _6893_ (.A(net323),
    .B(net243),
    .X(_3512_));
 sky130_fd_sc_hd__a31o_1 _6894_ (.A1(net458),
    .A2(net1885),
    .A3(net241),
    .B1(_3512_),
    .X(_1152_));
 sky130_fd_sc_hd__and2_1 _6895_ (.A(net325),
    .B(net244),
    .X(_3513_));
 sky130_fd_sc_hd__a31o_1 _6896_ (.A1(net461),
    .A2(net1666),
    .A3(_3503_),
    .B1(_3513_),
    .X(_1153_));
 sky130_fd_sc_hd__and2_1 _6897_ (.A(net324),
    .B(net243),
    .X(_3514_));
 sky130_fd_sc_hd__a31o_1 _6898_ (.A1(net459),
    .A2(net1758),
    .A3(net241),
    .B1(_3514_),
    .X(_1154_));
 sky130_fd_sc_hd__and2_1 _6899_ (.A(net322),
    .B(net244),
    .X(_3515_));
 sky130_fd_sc_hd__a31o_1 _6900_ (.A1(net453),
    .A2(net1703),
    .A3(net242),
    .B1(_3515_),
    .X(_1155_));
 sky130_fd_sc_hd__and2_1 _6901_ (.A(net319),
    .B(net243),
    .X(_3516_));
 sky130_fd_sc_hd__a31o_1 _6902_ (.A1(net459),
    .A2(net1920),
    .A3(net241),
    .B1(_3516_),
    .X(_1156_));
 sky130_fd_sc_hd__and2_1 _6903_ (.A(net321),
    .B(net244),
    .X(_3517_));
 sky130_fd_sc_hd__a31o_1 _6904_ (.A1(net454),
    .A2(net1760),
    .A3(net242),
    .B1(_3517_),
    .X(_1157_));
 sky130_fd_sc_hd__and2_1 _6905_ (.A(net320),
    .B(net243),
    .X(_3518_));
 sky130_fd_sc_hd__a31o_1 _6906_ (.A1(net452),
    .A2(net1836),
    .A3(net241),
    .B1(_3518_),
    .X(_1158_));
 sky130_fd_sc_hd__and2_1 _6907_ (.A(net318),
    .B(net243),
    .X(_3519_));
 sky130_fd_sc_hd__a31o_1 _6908_ (.A1(net458),
    .A2(net1848),
    .A3(net241),
    .B1(_3519_),
    .X(_1159_));
 sky130_fd_sc_hd__and2_1 _6909_ (.A(net342),
    .B(net244),
    .X(_3520_));
 sky130_fd_sc_hd__a31o_1 _6910_ (.A1(net453),
    .A2(net1696),
    .A3(net242),
    .B1(_3520_),
    .X(_1160_));
 sky130_fd_sc_hd__nor2_1 _6911_ (.A(_1381_),
    .B(net242),
    .Y(_3521_));
 sky130_fd_sc_hd__a31o_1 _6912_ (.A1(net444),
    .A2(net1544),
    .A3(net242),
    .B1(_3521_),
    .X(_1161_));
 sky130_fd_sc_hd__and2_1 _6913_ (.A(net341),
    .B(net243),
    .X(_3522_));
 sky130_fd_sc_hd__a31o_1 _6914_ (.A1(net460),
    .A2(net1828),
    .A3(net241),
    .B1(_3522_),
    .X(_1162_));
 sky130_fd_sc_hd__and2_1 _6915_ (.A(net343),
    .B(net244),
    .X(_3523_));
 sky130_fd_sc_hd__a31o_1 _6916_ (.A1(net450),
    .A2(net1658),
    .A3(net242),
    .B1(_3523_),
    .X(_1163_));
 sky130_fd_sc_hd__and2_1 _6917_ (.A(net338),
    .B(net244),
    .X(_3524_));
 sky130_fd_sc_hd__a31o_1 _6918_ (.A1(net445),
    .A2(net1778),
    .A3(net242),
    .B1(_3524_),
    .X(_1164_));
 sky130_fd_sc_hd__and2_1 _6919_ (.A(net340),
    .B(net244),
    .X(_3525_));
 sky130_fd_sc_hd__a31o_1 _6920_ (.A1(net447),
    .A2(net1748),
    .A3(net242),
    .B1(_3525_),
    .X(_1165_));
 sky130_fd_sc_hd__and2_1 _6921_ (.A(net339),
    .B(net243),
    .X(_3526_));
 sky130_fd_sc_hd__a31o_1 _6922_ (.A1(net455),
    .A2(net1939),
    .A3(net241),
    .B1(_3526_),
    .X(_1166_));
 sky130_fd_sc_hd__and2_1 _6923_ (.A(net337),
    .B(net244),
    .X(_3527_));
 sky130_fd_sc_hd__a31o_1 _6924_ (.A1(net446),
    .A2(net1783),
    .A3(net242),
    .B1(_3527_),
    .X(_1167_));
 sky130_fd_sc_hd__and2_1 _6925_ (.A(net334),
    .B(net243),
    .X(_3528_));
 sky130_fd_sc_hd__a31o_1 _6926_ (.A1(net461),
    .A2(net1810),
    .A3(net241),
    .B1(_3528_),
    .X(_1168_));
 sky130_fd_sc_hd__and2_1 _6927_ (.A(net336),
    .B(net244),
    .X(_3529_));
 sky130_fd_sc_hd__a31o_1 _6928_ (.A1(net446),
    .A2(net1793),
    .A3(net242),
    .B1(_3529_),
    .X(_1169_));
 sky130_fd_sc_hd__and2_1 _6929_ (.A(_1487_),
    .B(net244),
    .X(_3530_));
 sky130_fd_sc_hd__a31o_1 _6930_ (.A1(net446),
    .A2(net1711),
    .A3(net242),
    .B1(_3530_),
    .X(_1170_));
 sky130_fd_sc_hd__and2_1 _6931_ (.A(net333),
    .B(net244),
    .X(_3531_));
 sky130_fd_sc_hd__a31o_1 _6932_ (.A1(net454),
    .A2(net1602),
    .A3(net242),
    .B1(_3531_),
    .X(_1171_));
 sky130_fd_sc_hd__and2_1 _6933_ (.A(net346),
    .B(net244),
    .X(_3532_));
 sky130_fd_sc_hd__a31o_1 _6934_ (.A1(net447),
    .A2(net1791),
    .A3(net242),
    .B1(_3532_),
    .X(_1172_));
 sky130_fd_sc_hd__and2_1 _6935_ (.A(net344),
    .B(net244),
    .X(_3533_));
 sky130_fd_sc_hd__a31o_1 _6936_ (.A1(net445),
    .A2(net1822),
    .A3(net242),
    .B1(_3533_),
    .X(_1173_));
 sky130_fd_sc_hd__and2_1 _6937_ (.A(net345),
    .B(net243),
    .X(_3534_));
 sky130_fd_sc_hd__a31o_1 _6938_ (.A1(net461),
    .A2(net1856),
    .A3(net241),
    .B1(_3534_),
    .X(_1174_));
 sky130_fd_sc_hd__and2_1 _6939_ (.A(net368),
    .B(net244),
    .X(_3535_));
 sky130_fd_sc_hd__a31o_1 _6940_ (.A1(net448),
    .A2(net1528),
    .A3(net242),
    .B1(_3535_),
    .X(_1175_));
 sky130_fd_sc_hd__nor3_1 _6941_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2628_),
    .Y(_3536_));
 sky130_fd_sc_hd__or3_4 _6942_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2628_),
    .X(_3537_));
 sky130_fd_sc_hd__or3_1 _6943_ (.A(net472),
    .B(net2081),
    .C(net239),
    .X(_3538_));
 sky130_fd_sc_hd__o21a_1 _6944_ (.A1(_1564_),
    .A2(_3537_),
    .B1(_3538_),
    .X(_1176_));
 sky130_fd_sc_hd__and2_1 _6945_ (.A(_1548_),
    .B(net239),
    .X(_3539_));
 sky130_fd_sc_hd__a31o_1 _6946_ (.A1(net462),
    .A2(net1564),
    .A3(net237),
    .B1(_3539_),
    .X(_1177_));
 sky130_fd_sc_hd__and2_1 _6947_ (.A(_1535_),
    .B(net239),
    .X(_3540_));
 sky130_fd_sc_hd__a31o_1 _6948_ (.A1(net456),
    .A2(net1656),
    .A3(net237),
    .B1(_3540_),
    .X(_1178_));
 sky130_fd_sc_hd__and2_1 _6949_ (.A(net332),
    .B(net240),
    .X(_3541_));
 sky130_fd_sc_hd__a31o_1 _6950_ (.A1(net462),
    .A2(net1754),
    .A3(_3537_),
    .B1(_3541_),
    .X(_1179_));
 sky130_fd_sc_hd__and2_1 _6951_ (.A(_1584_),
    .B(net239),
    .X(_3542_));
 sky130_fd_sc_hd__a31o_1 _6952_ (.A1(net459),
    .A2(net1975),
    .A3(net237),
    .B1(_3542_),
    .X(_1180_));
 sky130_fd_sc_hd__or3b_1 _6953_ (.A(net470),
    .B(net239),
    .C_N(net2114),
    .X(_3543_));
 sky130_fd_sc_hd__o21ai_1 _6954_ (.A1(_1607_),
    .A2(net237),
    .B1(_3543_),
    .Y(_1181_));
 sky130_fd_sc_hd__and2_1 _6955_ (.A(_1596_),
    .B(net239),
    .X(_3544_));
 sky130_fd_sc_hd__a31o_1 _6956_ (.A1(net456),
    .A2(net1664),
    .A3(net237),
    .B1(_3544_),
    .X(_1182_));
 sky130_fd_sc_hd__and2_1 _6957_ (.A(net328),
    .B(net239),
    .X(_3545_));
 sky130_fd_sc_hd__a31o_1 _6958_ (.A1(net455),
    .A2(net1738),
    .A3(net237),
    .B1(_3545_),
    .X(_1183_));
 sky130_fd_sc_hd__and2_1 _6959_ (.A(_1644_),
    .B(net239),
    .X(_3546_));
 sky130_fd_sc_hd__a31o_1 _6960_ (.A1(net452),
    .A2(net1716),
    .A3(net237),
    .B1(_3546_),
    .X(_1184_));
 sky130_fd_sc_hd__and2_1 _6961_ (.A(_1624_),
    .B(net240),
    .X(_3547_));
 sky130_fd_sc_hd__a31o_1 _6962_ (.A1(net461),
    .A2(net1789),
    .A3(net237),
    .B1(_3547_),
    .X(_1185_));
 sky130_fd_sc_hd__and2_1 _6963_ (.A(_1633_),
    .B(net239),
    .X(_3548_));
 sky130_fd_sc_hd__a31o_1 _6964_ (.A1(net460),
    .A2(net1842),
    .A3(net237),
    .B1(_3548_),
    .X(_1186_));
 sky130_fd_sc_hd__and2_1 _6965_ (.A(_1655_),
    .B(net240),
    .X(_3549_));
 sky130_fd_sc_hd__a31o_1 _6966_ (.A1(net454),
    .A2(net1958),
    .A3(net238),
    .B1(_3549_),
    .X(_1187_));
 sky130_fd_sc_hd__and2_1 _6967_ (.A(_1690_),
    .B(net239),
    .X(_3550_));
 sky130_fd_sc_hd__a31o_1 _6968_ (.A1(net459),
    .A2(net1969),
    .A3(net237),
    .B1(_3550_),
    .X(_1188_));
 sky130_fd_sc_hd__and2_1 _6969_ (.A(_1667_),
    .B(net240),
    .X(_3551_));
 sky130_fd_sc_hd__a31o_1 _6970_ (.A1(net454),
    .A2(net1832),
    .A3(net238),
    .B1(_3551_),
    .X(_1189_));
 sky130_fd_sc_hd__and2_1 _6971_ (.A(net320),
    .B(net239),
    .X(_3552_));
 sky130_fd_sc_hd__a31o_1 _6972_ (.A1(net452),
    .A2(net1872),
    .A3(net237),
    .B1(_3552_),
    .X(_1190_));
 sky130_fd_sc_hd__and2_1 _6973_ (.A(_1702_),
    .B(net239),
    .X(_3553_));
 sky130_fd_sc_hd__a31o_1 _6974_ (.A1(net458),
    .A2(net1844),
    .A3(net237),
    .B1(_3553_),
    .X(_1191_));
 sky130_fd_sc_hd__and2_1 _6975_ (.A(_1407_),
    .B(net240),
    .X(_3554_));
 sky130_fd_sc_hd__a31o_1 _6976_ (.A1(net454),
    .A2(net1881),
    .A3(net238),
    .B1(_3554_),
    .X(_1192_));
 sky130_fd_sc_hd__nor2_1 _6977_ (.A(_1381_),
    .B(net238),
    .Y(_3555_));
 sky130_fd_sc_hd__a31o_1 _6978_ (.A1(net445),
    .A2(net1918),
    .A3(net238),
    .B1(_3555_),
    .X(_1193_));
 sky130_fd_sc_hd__and2_1 _6979_ (.A(_1420_),
    .B(net239),
    .X(_3556_));
 sky130_fd_sc_hd__a31o_1 _6980_ (.A1(net460),
    .A2(net1646),
    .A3(net237),
    .B1(_3556_),
    .X(_1194_));
 sky130_fd_sc_hd__and2_1 _6981_ (.A(_1396_),
    .B(net240),
    .X(_3557_));
 sky130_fd_sc_hd__a31o_1 _6982_ (.A1(net450),
    .A2(net1766),
    .A3(net238),
    .B1(_3557_),
    .X(_1195_));
 sky130_fd_sc_hd__and2_1 _6983_ (.A(net338),
    .B(net240),
    .X(_3558_));
 sky130_fd_sc_hd__a31o_1 _6984_ (.A1(net445),
    .A2(net1806),
    .A3(net238),
    .B1(_3558_),
    .X(_1196_));
 sky130_fd_sc_hd__and2_1 _6985_ (.A(_1432_),
    .B(net240),
    .X(_3559_));
 sky130_fd_sc_hd__a31o_1 _6986_ (.A1(net447),
    .A2(net1616),
    .A3(net238),
    .B1(_3559_),
    .X(_1197_));
 sky130_fd_sc_hd__and2_1 _6987_ (.A(net339),
    .B(net239),
    .X(_3560_));
 sky130_fd_sc_hd__a31o_1 _6988_ (.A1(net456),
    .A2(net1935),
    .A3(net237),
    .B1(_3560_),
    .X(_1198_));
 sky130_fd_sc_hd__and2_1 _6989_ (.A(net337),
    .B(net240),
    .X(_3561_));
 sky130_fd_sc_hd__a31o_1 _6990_ (.A1(net446),
    .A2(net1862),
    .A3(net238),
    .B1(_3561_),
    .X(_1199_));
 sky130_fd_sc_hd__and2_1 _6991_ (.A(_1498_),
    .B(net239),
    .X(_3562_));
 sky130_fd_sc_hd__a31o_1 _6992_ (.A1(net461),
    .A2(net1816),
    .A3(net237),
    .B1(_3562_),
    .X(_1200_));
 sky130_fd_sc_hd__and2_1 _6993_ (.A(_1475_),
    .B(net240),
    .X(_3563_));
 sky130_fd_sc_hd__a31o_1 _6994_ (.A1(net446),
    .A2(net1787),
    .A3(net238),
    .B1(_3563_),
    .X(_1201_));
 sky130_fd_sc_hd__and2_1 _6995_ (.A(net335),
    .B(net240),
    .X(_3564_));
 sky130_fd_sc_hd__a31o_1 _6996_ (.A1(net446),
    .A2(net1961),
    .A3(net238),
    .B1(_3564_),
    .X(_1202_));
 sky130_fd_sc_hd__and2_1 _6997_ (.A(_1510_),
    .B(net240),
    .X(_3565_));
 sky130_fd_sc_hd__a31o_1 _6998_ (.A1(net454),
    .A2(net1442),
    .A3(net238),
    .B1(_3565_),
    .X(_1203_));
 sky130_fd_sc_hd__and2_1 _6999_ (.A(_1343_),
    .B(net240),
    .X(_3566_));
 sky130_fd_sc_hd__a31o_1 _7000_ (.A1(net447),
    .A2(net1853),
    .A3(net238),
    .B1(_3566_),
    .X(_1204_));
 sky130_fd_sc_hd__and2_1 _7001_ (.A(_1366_),
    .B(net240),
    .X(_3567_));
 sky130_fd_sc_hd__a31o_1 _7002_ (.A1(net445),
    .A2(net1904),
    .A3(net238),
    .B1(_3567_),
    .X(_1205_));
 sky130_fd_sc_hd__and2_1 _7003_ (.A(_1355_),
    .B(net239),
    .X(_3568_));
 sky130_fd_sc_hd__a31o_1 _7004_ (.A1(net461),
    .A2(net1864),
    .A3(net237),
    .B1(_3568_),
    .X(_1206_));
 sky130_fd_sc_hd__and2_1 _7005_ (.A(_1316_),
    .B(net240),
    .X(_3569_));
 sky130_fd_sc_hd__a31o_1 _7006_ (.A1(net448),
    .A2(net1562),
    .A3(net238),
    .B1(_3569_),
    .X(_1207_));
 sky130_fd_sc_hd__nor2_1 _7007_ (.A(_2136_),
    .B(net162),
    .Y(_1208_));
 sky130_fd_sc_hd__or4_1 _7008_ (.A(net1990),
    .B(net1998),
    .C(net1698),
    .D(_2664_),
    .X(_3570_));
 sky130_fd_sc_hd__a21o_1 _7009_ (.A1(_0066_),
    .A2(_2663_),
    .B1(_2676_),
    .X(_3571_));
 sky130_fd_sc_hd__a2bb2o_1 _7010_ (.A1_N(net2091),
    .A2_N(_2672_),
    .B1(_2673_),
    .B2(_3571_),
    .X(_3572_));
 sky130_fd_sc_hd__a21boi_1 _7011_ (.A1(_2675_),
    .A2(_3572_),
    .B1_N(_2658_),
    .Y(_3573_));
 sky130_fd_sc_hd__o21ai_1 _7012_ (.A1(_2665_),
    .A2(_3573_),
    .B1(net2206),
    .Y(_3574_));
 sky130_fd_sc_hd__o211a_1 _7013_ (.A1(net2091),
    .A2(net2206),
    .B1(_3574_),
    .C1(_2646_),
    .X(_1209_));
 sky130_fd_sc_hd__a211o_1 _7014_ (.A1(net2091),
    .A2(net1698),
    .B1(_2669_),
    .C1(net1998),
    .X(_3575_));
 sky130_fd_sc_hd__a211o_1 _7015_ (.A1(_0067_),
    .A2(_2663_),
    .B1(_2671_),
    .C1(_2676_),
    .X(_3576_));
 sky130_fd_sc_hd__a21bo_1 _7016_ (.A1(_2670_),
    .A2(_3576_),
    .B1_N(_2672_),
    .X(_3577_));
 sky130_fd_sc_hd__a21bo_1 _7017_ (.A1(_3575_),
    .A2(_3577_),
    .B1_N(_2674_),
    .X(_3578_));
 sky130_fd_sc_hd__and3_1 _7018_ (.A(_2646_),
    .B(_2667_),
    .C(_3578_),
    .X(_1210_));
 sky130_fd_sc_hd__a22o_1 _7019_ (.A1(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ),
    .A2(_2671_),
    .B1(_2676_),
    .B2(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .X(_3579_));
 sky130_fd_sc_hd__a31o_1 _7020_ (.A1(_0064_),
    .A2(_2663_),
    .A3(_2677_),
    .B1(_3579_),
    .X(_3580_));
 sky130_fd_sc_hd__nand2_1 _7021_ (.A(_2654_),
    .B(_2660_),
    .Y(_3581_));
 sky130_fd_sc_hd__a32o_1 _7022_ (.A1(_2670_),
    .A2(_3580_),
    .A3(_3581_),
    .B1(_2668_),
    .B2(_2657_),
    .X(_3582_));
 sky130_fd_sc_hd__o211a_1 _7023_ (.A1(net2091),
    .A2(_2672_),
    .B1(_2675_),
    .C1(_3582_),
    .X(_3583_));
 sky130_fd_sc_hd__nor2_1 _7024_ (.A(_2666_),
    .B(_3583_),
    .Y(_3584_));
 sky130_fd_sc_hd__mux2_1 _7025_ (.A0(net2091),
    .A1(_3584_),
    .S(net2206),
    .X(_3585_));
 sky130_fd_sc_hd__nor2_1 _7026_ (.A(net162),
    .B(_3585_),
    .Y(_1211_));
 sky130_fd_sc_hd__nand2_1 _7027_ (.A(net1698),
    .B(_2656_),
    .Y(_3586_));
 sky130_fd_sc_hd__a221o_1 _7028_ (.A1(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .A2(_2655_),
    .B1(_2676_),
    .B2(net2205),
    .C1(_2671_),
    .X(_3587_));
 sky130_fd_sc_hd__a31o_1 _7029_ (.A1(_0065_),
    .A2(_2663_),
    .A3(_2677_),
    .B1(_3587_),
    .X(_3588_));
 sky130_fd_sc_hd__a21bo_1 _7030_ (.A1(_2669_),
    .A2(_3588_),
    .B1_N(_3575_),
    .X(_3589_));
 sky130_fd_sc_hd__a21oi_1 _7031_ (.A1(_3586_),
    .A2(_3589_),
    .B1(_2665_),
    .Y(_3590_));
 sky130_fd_sc_hd__mux2_1 _7032_ (.A0(net2091),
    .A1(_3590_),
    .S(net2206),
    .X(_3591_));
 sky130_fd_sc_hd__nor2_1 _7033_ (.A(net162),
    .B(_3591_),
    .Y(_1212_));
 sky130_fd_sc_hd__and2_1 _7034_ (.A(net462),
    .B(net1590),
    .X(_1213_));
 sky130_fd_sc_hd__and2_1 _7035_ (.A(net462),
    .B(net1552),
    .X(_1214_));
 sky130_fd_sc_hd__and2_1 _7036_ (.A(net456),
    .B(net1153),
    .X(_1215_));
 sky130_fd_sc_hd__and2_1 _7037_ (.A(net461),
    .B(net1289),
    .X(_1216_));
 sky130_fd_sc_hd__and2_1 _7038_ (.A(net459),
    .B(net1103),
    .X(_1217_));
 sky130_fd_sc_hd__and2_1 _7039_ (.A(net458),
    .B(net1403),
    .X(_1218_));
 sky130_fd_sc_hd__and2_1 _7040_ (.A(net456),
    .B(net1676),
    .X(_1219_));
 sky130_fd_sc_hd__and2_1 _7041_ (.A(net455),
    .B(net1209),
    .X(_1220_));
 sky130_fd_sc_hd__and2_1 _7042_ (.A(net458),
    .B(net1598),
    .X(_1221_));
 sky130_fd_sc_hd__and2_1 _7043_ (.A(net461),
    .B(net1426),
    .X(_1222_));
 sky130_fd_sc_hd__and2_1 _7044_ (.A(net460),
    .B(net1608),
    .X(_1223_));
 sky130_fd_sc_hd__and2_1 _7045_ (.A(net454),
    .B(net1707),
    .X(_1224_));
 sky130_fd_sc_hd__and2_1 _7046_ (.A(net459),
    .B(net1642),
    .X(_1225_));
 sky130_fd_sc_hd__and2_1 _7047_ (.A(net453),
    .B(net1377),
    .X(_1226_));
 sky130_fd_sc_hd__and2_1 _7048_ (.A(net452),
    .B(net1265),
    .X(_1227_));
 sky130_fd_sc_hd__and2_1 _7049_ (.A(net459),
    .B(net1682),
    .X(_1228_));
 sky130_fd_sc_hd__and2_1 _7050_ (.A(net453),
    .B(net1482),
    .X(_1229_));
 sky130_fd_sc_hd__and2_1 _7051_ (.A(net445),
    .B(net1630),
    .X(_1230_));
 sky130_fd_sc_hd__and2_1 _7052_ (.A(net460),
    .B(net1720),
    .X(_1231_));
 sky130_fd_sc_hd__and2_1 _7053_ (.A(net450),
    .B(net1341),
    .X(_1232_));
 sky130_fd_sc_hd__and2_1 _7054_ (.A(net445),
    .B(net1472),
    .X(_1233_));
 sky130_fd_sc_hd__and2_1 _7055_ (.A(net447),
    .B(net1087),
    .X(_1234_));
 sky130_fd_sc_hd__and2_1 _7056_ (.A(net456),
    .B(net1450),
    .X(_1235_));
 sky130_fd_sc_hd__and2_1 _7057_ (.A(net441),
    .B(net1594),
    .X(_1236_));
 sky130_fd_sc_hd__and2_1 _7058_ (.A(net461),
    .B(net1379),
    .X(_1237_));
 sky130_fd_sc_hd__and2_1 _7059_ (.A(net441),
    .B(net1600),
    .X(_1238_));
 sky130_fd_sc_hd__and2_1 _7060_ (.A(net446),
    .B(net1606),
    .X(_1239_));
 sky130_fd_sc_hd__and2_1 _7061_ (.A(net454),
    .B(net1053),
    .X(_1240_));
 sky130_fd_sc_hd__and2_1 _7062_ (.A(net447),
    .B(net1420),
    .X(_1241_));
 sky130_fd_sc_hd__and2_1 _7063_ (.A(net445),
    .B(net1538),
    .X(_1242_));
 sky130_fd_sc_hd__and2_1 _7064_ (.A(net461),
    .B(net1732),
    .X(_1243_));
 sky130_fd_sc_hd__and2_1 _7065_ (.A(net447),
    .B(net1512),
    .X(_1244_));
 sky130_fd_sc_hd__and3_1 _7066_ (.A(net1945),
    .B(net2085),
    .C(net276),
    .X(_1245_));
 sky130_fd_sc_hd__nand2_8 _7067_ (.A(net1945),
    .B(net2072),
    .Y(_3592_));
 sky130_fd_sc_hd__nand2_1 _7068_ (.A(net2091),
    .B(net2001),
    .Y(_3593_));
 sky130_fd_sc_hd__a21oi_1 _7069_ (.A1(_3592_),
    .A2(net2092),
    .B1(net162),
    .Y(_1246_));
 sky130_fd_sc_hd__nand2_1 _7070_ (.A(net2073),
    .B(net2001),
    .Y(_3594_));
 sky130_fd_sc_hd__a21oi_4 _7071_ (.A1(_3592_),
    .A2(_3594_),
    .B1(net162),
    .Y(_1247_));
 sky130_fd_sc_hd__nand2_1 _7072_ (.A(net1742),
    .B(net2001),
    .Y(_3595_));
 sky130_fd_sc_hd__a21oi_1 _7073_ (.A1(_3592_),
    .A2(net2002),
    .B1(net162),
    .Y(_1248_));
 sky130_fd_sc_hd__nand2_1 _7074_ (.A(net2116),
    .B(net2001),
    .Y(_3596_));
 sky130_fd_sc_hd__a21oi_1 _7075_ (.A1(_3592_),
    .A2(_3596_),
    .B1(net162),
    .Y(_1249_));
 sky130_fd_sc_hd__nand2_1 _7076_ (.A(net1972),
    .B(_2134_),
    .Y(_3597_));
 sky130_fd_sc_hd__a21oi_1 _7077_ (.A1(_3592_),
    .A2(net1973),
    .B1(net162),
    .Y(_1250_));
 sky130_fd_sc_hd__nand2_1 _7078_ (.A(net2018),
    .B(net2001),
    .Y(_3598_));
 sky130_fd_sc_hd__a21oi_1 _7079_ (.A1(_3592_),
    .A2(net2019),
    .B1(net162),
    .Y(_1251_));
 sky130_fd_sc_hd__nand2_1 _7080_ (.A(net2110),
    .B(net2001),
    .Y(_3599_));
 sky130_fd_sc_hd__a21oi_1 _7081_ (.A1(_3592_),
    .A2(net2111),
    .B1(net162),
    .Y(_1252_));
 sky130_fd_sc_hd__nand2_1 _7082_ (.A(net380),
    .B(net2001),
    .Y(_3600_));
 sky130_fd_sc_hd__a21oi_1 _7083_ (.A1(_3592_),
    .A2(net2113),
    .B1(net162),
    .Y(_1253_));
 sky130_fd_sc_hd__nand2_1 _7084_ (.A(net381),
    .B(net2001),
    .Y(_3601_));
 sky130_fd_sc_hd__a21oi_1 _7085_ (.A1(_3592_),
    .A2(net2099),
    .B1(net162),
    .Y(_1254_));
 sky130_fd_sc_hd__nand2_1 _7086_ (.A(net387),
    .B(net2001),
    .Y(_3602_));
 sky130_fd_sc_hd__a21oi_1 _7087_ (.A1(_3592_),
    .A2(net2097),
    .B1(net162),
    .Y(_1255_));
 sky130_fd_sc_hd__nand2_1 _7088_ (.A(net398),
    .B(net2001),
    .Y(_3603_));
 sky130_fd_sc_hd__a21oi_1 _7089_ (.A1(_3592_),
    .A2(net2090),
    .B1(net162),
    .Y(_1256_));
 sky130_fd_sc_hd__nand2_1 _7090_ (.A(net2126),
    .B(net2050),
    .Y(_3604_));
 sky130_fd_sc_hd__nand3_1 _7091_ (.A(net1945),
    .B(_2135_),
    .C(_2679_),
    .Y(_3605_));
 sky130_fd_sc_hd__a21oi_1 _7092_ (.A1(_3604_),
    .A2(net1946),
    .B1(net163),
    .Y(_1257_));
 sky130_fd_sc_hd__nand2_1 _7093_ (.A(net408),
    .B(_2680_),
    .Y(_3606_));
 sky130_fd_sc_hd__a21oi_1 _7094_ (.A1(net1946),
    .A2(_3606_),
    .B1(net163),
    .Y(_1258_));
 sky130_fd_sc_hd__nand2_1 _7095_ (.A(net414),
    .B(net2050),
    .Y(_3607_));
 sky130_fd_sc_hd__a21oi_1 _7096_ (.A1(net1946),
    .A2(_3607_),
    .B1(net163),
    .Y(_1259_));
 sky130_fd_sc_hd__nand2_1 _7097_ (.A(net419),
    .B(net2050),
    .Y(_3608_));
 sky130_fd_sc_hd__a21oi_1 _7098_ (.A1(net1946),
    .A2(_3608_),
    .B1(net163),
    .Y(_1260_));
 sky130_fd_sc_hd__nand2_1 _7099_ (.A(net428),
    .B(net2050),
    .Y(_3609_));
 sky130_fd_sc_hd__a21oi_1 _7100_ (.A1(net1946),
    .A2(net2051),
    .B1(net162),
    .Y(_1261_));
 sky130_fd_sc_hd__nand2_1 _7101_ (.A(net1990),
    .B(_2680_),
    .Y(_3610_));
 sky130_fd_sc_hd__a21oi_1 _7102_ (.A1(net1946),
    .A2(net1991),
    .B1(net163),
    .Y(_1262_));
 sky130_fd_sc_hd__nand2_1 _7103_ (.A(net1998),
    .B(_2680_),
    .Y(_3611_));
 sky130_fd_sc_hd__a21oi_1 _7104_ (.A1(net1946),
    .A2(net1999),
    .B1(net163),
    .Y(_1263_));
 sky130_fd_sc_hd__nand2_1 _7105_ (.A(net1698),
    .B(_2680_),
    .Y(_3612_));
 sky130_fd_sc_hd__a21oi_1 _7106_ (.A1(_3605_),
    .A2(net1699),
    .B1(net163),
    .Y(_1264_));
 sky130_fd_sc_hd__nor2_1 _7107_ (.A(_2660_),
    .B(net1946),
    .Y(_3613_));
 sky130_fd_sc_hd__a32o_1 _7108_ (.A1(net398),
    .A2(net2048),
    .A3(_2132_),
    .B1(_2660_),
    .B2(net877),
    .X(_3614_));
 sky130_fd_sc_hd__o21a_1 _7109_ (.A1(_3613_),
    .A2(_3614_),
    .B1(_2646_),
    .X(_1265_));
 sky130_fd_sc_hd__and3_1 _7110_ (.A(net2091),
    .B(net2072),
    .C(_2646_),
    .X(_1266_));
 sky130_fd_sc_hd__and3_1 _7111_ (.A(net2073),
    .B(net2072),
    .C(_2646_),
    .X(_1267_));
 sky130_fd_sc_hd__and3_1 _7112_ (.A(net1742),
    .B(_2135_),
    .C(_2646_),
    .X(_1268_));
 sky130_fd_sc_hd__and3_1 _7113_ (.A(net2116),
    .B(net2072),
    .C(_2646_),
    .X(_1269_));
 sky130_fd_sc_hd__and3_1 _7114_ (.A(net1972),
    .B(net2072),
    .C(_2646_),
    .X(_1270_));
 sky130_fd_sc_hd__and3_1 _7115_ (.A(net2018),
    .B(net2072),
    .C(_2646_),
    .X(_1271_));
 sky130_fd_sc_hd__nor2_1 _7116_ (.A(_2659_),
    .B(_2680_),
    .Y(_3615_));
 sky130_fd_sc_hd__o21ai_2 _7117_ (.A1(_2134_),
    .A2(_2659_),
    .B1(_2679_),
    .Y(_3616_));
 sky130_fd_sc_hd__a22o_1 _7118_ (.A1(net2131),
    .A2(_2659_),
    .B1(_3616_),
    .B2(net2110),
    .X(_3617_));
 sky130_fd_sc_hd__and3_1 _7119_ (.A(net175),
    .B(net277),
    .C(_3617_),
    .X(_1272_));
 sky130_fd_sc_hd__a22o_1 _7120_ (.A1(net2107),
    .A2(_2659_),
    .B1(_3616_),
    .B2(net380),
    .X(_3618_));
 sky130_fd_sc_hd__and3_1 _7121_ (.A(net176),
    .B(net280),
    .C(_3618_),
    .X(_1273_));
 sky130_fd_sc_hd__a22o_1 _7122_ (.A1(net2153),
    .A2(_2659_),
    .B1(_3616_),
    .B2(net382),
    .X(_3619_));
 sky130_fd_sc_hd__and3_1 _7123_ (.A(net176),
    .B(net277),
    .C(_3619_),
    .X(_1274_));
 sky130_fd_sc_hd__a22o_1 _7124_ (.A1(net2151),
    .A2(_2659_),
    .B1(_3616_),
    .B2(net389),
    .X(_3620_));
 sky130_fd_sc_hd__and3_1 _7125_ (.A(net176),
    .B(net277),
    .C(_3620_),
    .X(_1275_));
 sky130_fd_sc_hd__a32o_1 _7126_ (.A1(net877),
    .A2(_1277_),
    .A3(_2659_),
    .B1(_3615_),
    .B2(net400),
    .X(_3621_));
 sky130_fd_sc_hd__and3_1 _7127_ (.A(net175),
    .B(net277),
    .C(_3621_),
    .X(_1276_));
 sky130_fd_sc_hd__o31a_1 _7128_ (.A1(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .A2(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .A3(_2137_),
    .B1(_2136_),
    .X(_3624_));
 sky130_fd_sc_hd__o31a_1 _7129_ (.A1(net2202),
    .A2(net2309),
    .A3(_2137_),
    .B1(_2136_),
    .X(_3625_));
 sky130_fd_sc_hd__o31a_1 _7130_ (.A1(net2124),
    .A2(net2071),
    .A3(_2137_),
    .B1(_2136_),
    .X(_3626_));
 sky130_fd_sc_hd__o31a_1 _7131_ (.A1(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .A2(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .A3(_2137_),
    .B1(_2136_),
    .X(_3622_));
 sky130_fd_sc_hd__inv_2 _7132_ (.A(net470),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _7133_ (.A(net470),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _7134_ (.A(net468),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _7135_ (.A(net468),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _7136_ (.A(net470),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _7137_ (.A(net470),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _7138_ (.A(net470),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _7139_ (.A(net468),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _7140_ (.A(net468),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _7141_ (.A(net470),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _7142_ (.A(net469),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _7143_ (.A(net468),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _7144_ (.A(net470),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _7145_ (.A(net468),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _7146_ (.A(net469),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _7147_ (.A(net470),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _7148_ (.A(net469),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _7149_ (.A(net464),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _7150_ (.A(net464),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _7151_ (.A(net465),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _7152_ (.A(net464),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _7153_ (.A(net465),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _7154_ (.A(net464),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _7155_ (.A(net465),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _7156_ (.A(net464),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _7157_ (.A(net464),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _7158_ (.A(net466),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _7159_ (.A(net464),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _7160_ (.A(net464),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _7161__2 (.A(clknet_leaf_38_clk),
    .Y(net481));
 sky130_fd_sc_hd__inv_2 _7162__3 (.A(clknet_leaf_40_clk),
    .Y(net482));
 sky130_fd_sc_hd__inv_2 _7163__4 (.A(clknet_leaf_33_clk),
    .Y(net483));
 sky130_fd_sc_hd__inv_2 _7164__5 (.A(clknet_leaf_27_clk),
    .Y(net484));
 sky130_fd_sc_hd__inv_2 _7165__6 (.A(clknet_leaf_26_clk),
    .Y(net485));
 sky130_fd_sc_hd__inv_2 _7166__7 (.A(clknet_leaf_41_clk),
    .Y(net486));
 sky130_fd_sc_hd__inv_2 _7167__8 (.A(clknet_leaf_48_clk),
    .Y(net487));
 sky130_fd_sc_hd__inv_2 _7168__9 (.A(clknet_leaf_22_clk),
    .Y(net488));
 sky130_fd_sc_hd__inv_2 _7169__10 (.A(clknet_leaf_33_clk),
    .Y(net489));
 sky130_fd_sc_hd__inv_2 _7170__11 (.A(clknet_leaf_25_clk),
    .Y(net490));
 sky130_fd_sc_hd__inv_2 _7171__12 (.A(clknet_leaf_56_clk),
    .Y(net491));
 sky130_fd_sc_hd__inv_2 _7172__13 (.A(clknet_leaf_12_clk),
    .Y(net492));
 sky130_fd_sc_hd__inv_2 _7173__14 (.A(clknet_leaf_43_clk),
    .Y(net493));
 sky130_fd_sc_hd__inv_2 _7174__15 (.A(clknet_leaf_21_clk),
    .Y(net494));
 sky130_fd_sc_hd__inv_2 _7175__16 (.A(clknet_leaf_26_clk),
    .Y(net495));
 sky130_fd_sc_hd__inv_2 _7176__17 (.A(clknet_leaf_45_clk),
    .Y(net496));
 sky130_fd_sc_hd__inv_2 _7177__18 (.A(clknet_leaf_54_clk),
    .Y(net497));
 sky130_fd_sc_hd__inv_2 _7178__19 (.A(clknet_leaf_24_clk),
    .Y(net498));
 sky130_fd_sc_hd__inv_2 _7179__20 (.A(clknet_leaf_51_clk),
    .Y(net499));
 sky130_fd_sc_hd__inv_2 _7180__21 (.A(clknet_leaf_55_clk),
    .Y(net500));
 sky130_fd_sc_hd__inv_2 _7181__22 (.A(clknet_leaf_60_clk),
    .Y(net501));
 sky130_fd_sc_hd__inv_2 _7182__23 (.A(clknet_leaf_46_clk),
    .Y(net502));
 sky130_fd_sc_hd__inv_2 _7183__24 (.A(clknet_leaf_62_clk),
    .Y(net503));
 sky130_fd_sc_hd__inv_2 _7184__25 (.A(clknet_leaf_31_clk),
    .Y(net504));
 sky130_fd_sc_hd__inv_2 _7185__26 (.A(clknet_leaf_62_clk),
    .Y(net505));
 sky130_fd_sc_hd__inv_2 _7186__27 (.A(clknet_leaf_61_clk),
    .Y(net506));
 sky130_fd_sc_hd__inv_2 _7187__28 (.A(clknet_leaf_43_clk),
    .Y(net507));
 sky130_fd_sc_hd__inv_2 _7188__29 (.A(clknet_leaf_55_clk),
    .Y(net508));
 sky130_fd_sc_hd__inv_2 _7189__30 (.A(clknet_leaf_75_clk),
    .Y(net509));
 sky130_fd_sc_hd__inv_2 _7190__31 (.A(clknet_leaf_29_clk),
    .Y(net510));
 sky130_fd_sc_hd__inv_2 _7191__32 (.A(clknet_leaf_58_clk),
    .Y(net511));
 sky130_fd_sc_hd__inv_2 _7192__33 (.A(clknet_leaf_38_clk),
    .Y(net512));
 sky130_fd_sc_hd__inv_2 _7193__34 (.A(clknet_leaf_38_clk),
    .Y(net513));
 sky130_fd_sc_hd__inv_2 _7194__35 (.A(clknet_leaf_39_clk),
    .Y(net514));
 sky130_fd_sc_hd__inv_2 _7195__36 (.A(clknet_leaf_33_clk),
    .Y(net515));
 sky130_fd_sc_hd__inv_2 _7196__37 (.A(clknet_leaf_12_clk),
    .Y(net516));
 sky130_fd_sc_hd__inv_2 _7197__38 (.A(clknet_leaf_13_clk),
    .Y(net517));
 sky130_fd_sc_hd__inv_2 _7198__39 (.A(clknet_leaf_40_clk),
    .Y(net518));
 sky130_fd_sc_hd__inv_2 _7199__40 (.A(clknet_leaf_23_clk),
    .Y(net519));
 sky130_fd_sc_hd__inv_2 _7200__41 (.A(clknet_leaf_22_clk),
    .Y(net520));
 sky130_fd_sc_hd__inv_2 _7201__42 (.A(clknet_leaf_33_clk),
    .Y(net521));
 sky130_fd_sc_hd__inv_2 _7202__43 (.A(clknet_leaf_24_clk),
    .Y(net522));
 sky130_fd_sc_hd__inv_2 _7203__44 (.A(clknet_leaf_57_clk),
    .Y(net523));
 sky130_fd_sc_hd__inv_2 _7204__45 (.A(clknet_leaf_12_clk),
    .Y(net524));
 sky130_fd_sc_hd__inv_2 _7205__46 (.A(clknet_leaf_44_clk),
    .Y(net525));
 sky130_fd_sc_hd__inv_2 _7206__47 (.A(clknet_leaf_21_clk),
    .Y(net526));
 sky130_fd_sc_hd__inv_2 _7207__48 (.A(clknet_leaf_26_clk),
    .Y(net527));
 sky130_fd_sc_hd__inv_2 _7208__49 (.A(clknet_leaf_49_clk),
    .Y(net528));
 sky130_fd_sc_hd__inv_2 _7209__50 (.A(clknet_leaf_54_clk),
    .Y(net529));
 sky130_fd_sc_hd__inv_2 _7210__51 (.A(clknet_leaf_32_clk),
    .Y(net530));
 sky130_fd_sc_hd__inv_2 _7211__52 (.A(clknet_leaf_50_clk),
    .Y(net531));
 sky130_fd_sc_hd__inv_2 _7212__53 (.A(clknet_leaf_55_clk),
    .Y(net532));
 sky130_fd_sc_hd__inv_2 _7213__54 (.A(clknet_leaf_58_clk),
    .Y(net533));
 sky130_fd_sc_hd__inv_2 _7214__55 (.A(clknet_leaf_46_clk),
    .Y(net534));
 sky130_fd_sc_hd__inv_2 _7215__56 (.A(clknet_leaf_61_clk),
    .Y(net535));
 sky130_fd_sc_hd__inv_2 _7216__57 (.A(clknet_leaf_31_clk),
    .Y(net536));
 sky130_fd_sc_hd__inv_2 _7217__58 (.A(clknet_leaf_62_clk),
    .Y(net537));
 sky130_fd_sc_hd__inv_2 _7218__59 (.A(clknet_leaf_62_clk),
    .Y(net538));
 sky130_fd_sc_hd__inv_2 _7219__60 (.A(clknet_leaf_44_clk),
    .Y(net539));
 sky130_fd_sc_hd__inv_2 _7220__61 (.A(clknet_leaf_75_clk),
    .Y(net540));
 sky130_fd_sc_hd__inv_2 _7221__62 (.A(clknet_leaf_74_clk),
    .Y(net541));
 sky130_fd_sc_hd__inv_2 _7222__63 (.A(clknet_leaf_31_clk),
    .Y(net542));
 sky130_fd_sc_hd__inv_2 _7223__64 (.A(clknet_leaf_58_clk),
    .Y(net543));
 sky130_fd_sc_hd__inv_2 _7224_ (.A(net466),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _7225_ (.A(net470),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _7226_ (.A(net470),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _7227_ (.A(net469),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _7228_ (.A(net470),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _7229_ (.A(net470),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _7230_ (.A(net470),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _7231_ (.A(net63),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _7232_ (.A(net469),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _7233_ (.A(net468),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _7234_ (.A(net469),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _7235_ (.A(net468),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _7236_ (.A(net468),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _7237_ (.A(net468),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _7238_ (.A(net469),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _7239_ (.A(net469),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _7240_ (.A(net469),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _7241_ (.A(net469),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _7242_ (.A(net467),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _7243_ (.A(net465),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _7244_ (.A(net465),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _7245_ (.A(net465),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _7246_ (.A(net465),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _7247_ (.A(net464),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _7248_ (.A(net465),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _7249_ (.A(net464),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _7250_ (.A(net464),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _7251_ (.A(net464),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _7252_ (.A(net464),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _7253_ (.A(net464),
    .Y(_0192_));
 sky130_fd_sc_hd__dfxtp_1 _7254_ (.CLK(clknet_leaf_73_clk),
    .D(net745),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7255_ (.CLK(clknet_leaf_17_clk),
    .D(net1995),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7256_ (.CLK(clknet_leaf_18_clk),
    .D(net2120),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7257_ (.CLK(clknet_leaf_7_clk),
    .D(net2117),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7258_ (.CLK(clknet_leaf_19_clk),
    .D(net2035),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7259_ (.CLK(clknet_leaf_7_clk),
    .D(net1417),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7260_ (.CLK(clknet_3_4_0_clk),
    .D(net2242),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7261_ (.CLK(clknet_leaf_15_clk),
    .D(net2069),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7262_ (.CLK(clknet_leaf_2_clk),
    .D(net2088),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7263_ (.CLK(clknet_leaf_6_clk),
    .D(net2011),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7264_ (.CLK(clknet_leaf_11_clk),
    .D(net1780),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7265_ (.CLK(clknet_leaf_48_clk),
    .D(net809),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7266_ (.CLK(clknet_leaf_19_clk),
    .D(net2046),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7267_ (.CLK(clknet_leaf_15_clk),
    .D(net1901),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7268_ (.CLK(clknet_leaf_51_clk),
    .D(net2123),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7269_ (.CLK(clknet_leaf_48_clk),
    .D(net1944),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7270_ (.CLK(clknet_leaf_13_clk),
    .D(net1943),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7271_ (.CLK(clknet_leaf_53_clk),
    .D(net1797),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7272_ (.CLK(clknet_leaf_71_clk),
    .D(net779),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7273_ (.CLK(clknet_leaf_63_clk),
    .D(net2095),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7274_ (.CLK(clknet_leaf_63_clk),
    .D(net2119),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7275_ (.CLK(clknet_leaf_71_clk),
    .D(net929),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7276_ (.CLK(clknet_leaf_68_clk),
    .D(net1997),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7277_ (.CLK(clknet_leaf_67_clk),
    .D(net796),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7278_ (.CLK(clknet_leaf_68_clk),
    .D(net1713),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7279_ (.CLK(clknet_leaf_70_clk),
    .D(net2179),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7280_ (.CLK(clknet_leaf_71_clk),
    .D(net1850),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7281_ (.CLK(clknet_leaf_72_clk),
    .D(net1960),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7282_ (.CLK(clknet_leaf_70_clk),
    .D(net2012),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7283_ (.CLK(clknet_leaf_67_clk),
    .D(net2106),
    .Q(\U_DATAPATH.U_IF_ID.i_pc_IF[31] ));
 sky130_fd_sc_hd__dfxtp_4 _7284_ (.CLK(clknet_leaf_77_clk),
    .D(net635),
    .Q(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__dfxtp_4 _7285_ (.CLK(clknet_leaf_4_clk),
    .D(net672),
    .Q(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7286_ (.CLK(clknet_leaf_73_clk),
    .D(_0195_),
    .RESET_B(net437),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_4 _7287_ (.CLK(clknet_leaf_17_clk),
    .D(_0196_),
    .RESET_B(_0070_),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_4 _7288_ (.CLK(clknet_leaf_17_clk),
    .D(_0197_),
    .RESET_B(_0071_),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_4 _7289_ (.CLK(clknet_leaf_7_clk),
    .D(_0198_),
    .RESET_B(_0072_),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_4 _7290_ (.CLK(clknet_leaf_6_clk),
    .D(_0199_),
    .RESET_B(_0073_),
    .Q(net126));
 sky130_fd_sc_hd__dfrtp_4 _7291_ (.CLK(clknet_leaf_16_clk),
    .D(_0200_),
    .RESET_B(_0074_),
    .Q(net127));
 sky130_fd_sc_hd__dfrtp_4 _7292_ (.CLK(clknet_leaf_16_clk),
    .D(_0201_),
    .RESET_B(_0075_),
    .Q(net128));
 sky130_fd_sc_hd__dfrtp_4 _7293_ (.CLK(clknet_leaf_15_clk),
    .D(_0202_),
    .RESET_B(_0076_),
    .Q(net129));
 sky130_fd_sc_hd__dfrtp_4 _7294_ (.CLK(clknet_leaf_2_clk),
    .D(_0203_),
    .RESET_B(_0077_),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_4 _7295_ (.CLK(clknet_leaf_6_clk),
    .D(_0204_),
    .RESET_B(_0078_),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_4 _7296_ (.CLK(clknet_leaf_11_clk),
    .D(_0205_),
    .RESET_B(_0079_),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_4 _7297_ (.CLK(clknet_leaf_50_clk),
    .D(_0206_),
    .RESET_B(_0080_),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_4 _7298_ (.CLK(clknet_leaf_5_clk),
    .D(_0207_),
    .RESET_B(_0081_),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_4 _7299_ (.CLK(clknet_leaf_15_clk),
    .D(_0208_),
    .RESET_B(_0082_),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_4 _7300_ (.CLK(clknet_leaf_21_clk),
    .D(_0209_),
    .RESET_B(_0083_),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_4 _7301_ (.CLK(clknet_leaf_48_clk),
    .D(_0210_),
    .RESET_B(_0084_),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_4 _7302_ (.CLK(clknet_leaf_13_clk),
    .D(_0211_),
    .RESET_B(_0085_),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_4 _7303_ (.CLK(clknet_leaf_53_clk),
    .D(_0212_),
    .RESET_B(_0086_),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_1 _7304_ (.CLK(clknet_leaf_71_clk),
    .D(_0213_),
    .RESET_B(_0087_),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_4 _7305_ (.CLK(clknet_leaf_63_clk),
    .D(_0214_),
    .RESET_B(_0088_),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_4 _7306_ (.CLK(clknet_leaf_63_clk),
    .D(_0215_),
    .RESET_B(_0089_),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_4 _7307_ (.CLK(clknet_leaf_67_clk),
    .D(_0216_),
    .RESET_B(_0090_),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_4 _7308_ (.CLK(clknet_leaf_68_clk),
    .D(_0217_),
    .RESET_B(_0091_),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_2 _7309_ (.CLK(clknet_leaf_67_clk),
    .D(_0218_),
    .RESET_B(_0092_),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_4 _7310_ (.CLK(clknet_leaf_68_clk),
    .D(_0219_),
    .RESET_B(_0093_),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_4 _7311_ (.CLK(clknet_leaf_68_clk),
    .D(_0220_),
    .RESET_B(_0094_),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_4 _7312_ (.CLK(clknet_leaf_71_clk),
    .D(_0221_),
    .RESET_B(_0095_),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_4 _7313_ (.CLK(clknet_leaf_72_clk),
    .D(_0222_),
    .RESET_B(_0096_),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_4 _7314_ (.CLK(clknet_leaf_70_clk),
    .D(_0223_),
    .RESET_B(_0097_),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_4 _7315_ (.CLK(clknet_leaf_70_clk),
    .D(_0224_),
    .RESET_B(_0098_),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_1 _7316_ (.CLK(clknet_leaf_73_clk),
    .D(net2101),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7317_ (.CLK(clknet_leaf_16_clk),
    .D(_0226_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7318_ (.CLK(clknet_leaf_16_clk),
    .D(_0227_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7319_ (.CLK(clknet_leaf_7_clk),
    .D(_0228_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7320_ (.CLK(clknet_leaf_17_clk),
    .D(_0229_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7321_ (.CLK(clknet_leaf_15_clk),
    .D(_0230_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7322_ (.CLK(clknet_leaf_16_clk),
    .D(_0231_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7323_ (.CLK(clknet_leaf_15_clk),
    .D(_0232_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7324_ (.CLK(clknet_leaf_6_clk),
    .D(_0233_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7325_ (.CLK(clknet_leaf_6_clk),
    .D(_0234_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7326_ (.CLK(clknet_leaf_15_clk),
    .D(_0235_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7327_ (.CLK(clknet_leaf_4_clk),
    .D(_0236_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7328_ (.CLK(clknet_leaf_6_clk),
    .D(_0237_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7329_ (.CLK(clknet_leaf_6_clk),
    .D(_0238_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7330_ (.CLK(clknet_leaf_48_clk),
    .D(_0239_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7331_ (.CLK(clknet_leaf_20_clk),
    .D(_0240_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7332_ (.CLK(clknet_leaf_47_clk),
    .D(_0241_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7333_ (.CLK(clknet_leaf_53_clk),
    .D(_0242_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7334_ (.CLK(clknet_leaf_75_clk),
    .D(_0243_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7335_ (.CLK(clknet_leaf_64_clk),
    .D(net1875),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7336_ (.CLK(clknet_leaf_69_clk),
    .D(_0245_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7337_ (.CLK(clknet_leaf_64_clk),
    .D(_0246_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7338_ (.CLK(clknet_leaf_68_clk),
    .D(_0247_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7339_ (.CLK(clknet_leaf_67_clk),
    .D(_0248_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7340_ (.CLK(clknet_leaf_68_clk),
    .D(_0249_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7341_ (.CLK(clknet_leaf_68_clk),
    .D(_0250_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7342_ (.CLK(clknet_leaf_72_clk),
    .D(net1955),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7343_ (.CLK(clknet_leaf_71_clk),
    .D(_0252_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7344_ (.CLK(clknet_leaf_72_clk),
    .D(net1888),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7345_ (.CLK(clknet_leaf_71_clk),
    .D(_0254_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7346_ (.CLK(clknet_leaf_3_clk),
    .D(_0255_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7347_ (.CLK(clknet_leaf_2_clk),
    .D(_0256_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7348_ (.CLK(clknet_leaf_2_clk),
    .D(_0257_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7349_ (.CLK(clknet_leaf_2_clk),
    .D(_0258_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7350_ (.CLK(clknet_leaf_2_clk),
    .D(_0259_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7351_ (.CLK(clknet_leaf_11_clk),
    .D(_0260_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7352_ (.CLK(clknet_leaf_6_clk),
    .D(_0261_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7353_ (.CLK(clknet_leaf_37_clk),
    .D(_0262_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7354_ (.CLK(clknet_leaf_11_clk),
    .D(_0263_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7355_ (.CLK(clknet_leaf_1_clk),
    .D(_0264_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[11] ));
 sky130_fd_sc_hd__dfxtp_2 _7356_ (.CLK(clknet_leaf_80_clk),
    .D(_0265_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7357_ (.CLK(clknet_leaf_11_clk),
    .D(_0266_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7358_ (.CLK(clknet_leaf_12_clk),
    .D(_0267_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__dfxtp_4 _7359_ (.CLK(clknet_leaf_12_clk),
    .D(_0268_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__dfxtp_4 _7360_ (.CLK(clknet_leaf_60_clk),
    .D(_0269_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7361_ (.CLK(clknet_leaf_71_clk),
    .D(_0270_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7362_ (.CLK(clknet_leaf_73_clk),
    .D(_0271_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7363_ (.CLK(clknet_leaf_43_clk),
    .D(_0272_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7364_ (.CLK(clknet_leaf_35_clk),
    .D(_0273_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7365_ (.CLK(clknet_leaf_61_clk),
    .D(_0274_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7366_ (.CLK(clknet_leaf_36_clk),
    .D(_0275_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ));
 sky130_fd_sc_hd__dfxtp_4 _7367_ (.CLK(clknet_leaf_65_clk),
    .D(_0276_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7368_ (.CLK(clknet_leaf_41_clk),
    .D(_0277_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7369_ (.CLK(clknet_leaf_1_clk),
    .D(_0278_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7370_ (.CLK(clknet_leaf_73_clk),
    .D(_0279_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7371_ (.CLK(clknet_leaf_59_clk),
    .D(_0280_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7372_ (.CLK(clknet_leaf_82_clk),
    .D(_0281_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7373_ (.CLK(clknet_leaf_28_clk),
    .D(_0282_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7374_ (.CLK(clknet_leaf_66_clk),
    .D(_0283_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ));
 sky130_fd_sc_hd__dfxtp_1 _7375_ (.CLK(clknet_leaf_1_clk),
    .D(_0284_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7376_ (.CLK(clknet_leaf_73_clk),
    .D(net922),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7377_ (.CLK(clknet_leaf_18_clk),
    .D(net712),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7378_ (.CLK(clknet_leaf_18_clk),
    .D(net881),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7379_ (.CLK(clknet_leaf_7_clk),
    .D(net866),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7380_ (.CLK(clknet_leaf_19_clk),
    .D(net851),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7381_ (.CLK(clknet_leaf_7_clk),
    .D(net825),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7382_ (.CLK(clknet_leaf_7_clk),
    .D(net545),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7383_ (.CLK(clknet_leaf_15_clk),
    .D(net959),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7384_ (.CLK(clknet_leaf_2_clk),
    .D(net976),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7385_ (.CLK(clknet_leaf_6_clk),
    .D(net845),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7386_ (.CLK(clknet_leaf_11_clk),
    .D(net827),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7387_ (.CLK(clknet_leaf_49_clk),
    .D(net783),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7388_ (.CLK(clknet_leaf_19_clk),
    .D(net831),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7389_ (.CLK(clknet_leaf_15_clk),
    .D(net891),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7390_ (.CLK(clknet_leaf_51_clk),
    .D(net817),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7391_ (.CLK(clknet_leaf_48_clk),
    .D(net972),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7392_ (.CLK(clknet_leaf_13_clk),
    .D(net859),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7393_ (.CLK(clknet_leaf_57_clk),
    .D(net647),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7394_ (.CLK(clknet_leaf_71_clk),
    .D(net889),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7395_ (.CLK(clknet_leaf_63_clk),
    .D(net862),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7396_ (.CLK(clknet_leaf_63_clk),
    .D(net855),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7397_ (.CLK(clknet_leaf_67_clk),
    .D(net777),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7398_ (.CLK(clknet_leaf_64_clk),
    .D(net761),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7399_ (.CLK(clknet_leaf_67_clk),
    .D(net947),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7400_ (.CLK(clknet_leaf_68_clk),
    .D(net897),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7401_ (.CLK(clknet_leaf_70_clk),
    .D(net829),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7402_ (.CLK(clknet_leaf_71_clk),
    .D(net847),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7403_ (.CLK(clknet_leaf_72_clk),
    .D(net1012),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7404_ (.CLK(clknet_leaf_70_clk),
    .D(net837),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7405_ (.CLK(clknet_leaf_67_clk),
    .D(net819),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7406_ (.CLK(clknet_leaf_38_clk),
    .D(net937),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7407_ (.CLK(clknet_leaf_35_clk),
    .D(net1026),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7408_ (.CLK(clknet_leaf_38_clk),
    .D(net996),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7409_ (.CLK(clknet_leaf_38_clk),
    .D(net1725),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7410_ (.CLK(clknet_leaf_27_clk),
    .D(net1074),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7411_ (.CLK(clknet_leaf_25_clk),
    .D(net1489),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7412_ (.CLK(clknet_leaf_39_clk),
    .D(net1116),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7413_ (.CLK(clknet_leaf_23_clk),
    .D(net1463),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7414_ (.CLK(clknet_leaf_22_clk),
    .D(net1114),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7415_ (.CLK(clknet_leaf_33_clk),
    .D(net1459),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7416_ (.CLK(clknet_leaf_24_clk),
    .D(net1166),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7417_ (.CLK(clknet_leaf_57_clk),
    .D(net1431),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7418_ (.CLK(clknet_leaf_31_clk),
    .D(net1573),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7419_ (.CLK(clknet_leaf_44_clk),
    .D(net1673),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7420_ (.CLK(clknet_leaf_21_clk),
    .D(net1715),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7421_ (.CLK(clknet_leaf_27_clk),
    .D(net1216),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7422_ (.CLK(clknet_leaf_48_clk),
    .D(net1481),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7423_ (.CLK(clknet_leaf_54_clk),
    .D(net1100),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7424_ (.CLK(clknet_leaf_31_clk),
    .D(net1352),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7425_ (.CLK(clknet_leaf_50_clk),
    .D(net1120),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7426_ (.CLK(clknet_leaf_56_clk),
    .D(net1517),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7427_ (.CLK(clknet_leaf_57_clk),
    .D(net1134),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7428_ (.CLK(clknet_leaf_46_clk),
    .D(net1597),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7429_ (.CLK(clknet_leaf_58_clk),
    .D(net1168),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7430_ (.CLK(clknet_leaf_31_clk),
    .D(net1497),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7431_ (.CLK(clknet_leaf_56_clk),
    .D(net1547),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7432_ (.CLK(clknet_leaf_58_clk),
    .D(net1130),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7433_ (.CLK(clknet_leaf_44_clk),
    .D(net1465),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7434_ (.CLK(clknet_leaf_57_clk),
    .D(net1094),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7435_ (.CLK(clknet_leaf_54_clk),
    .D(net1613),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7436_ (.CLK(clknet_leaf_31_clk),
    .D(net1737),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7437_ (.CLK(clknet_leaf_58_clk),
    .D(net966),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7438_ (.CLK(clknet_leaf_38_clk),
    .D(net1521),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7439_ (.CLK(clknet_leaf_33_clk),
    .D(net1048),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7440_ (.CLK(clknet_leaf_39_clk),
    .D(net1382),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7441_ (.CLK(clknet_leaf_33_clk),
    .D(net870),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7442_ (.CLK(clknet_leaf_28_clk),
    .D(net1102),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7443_ (.CLK(clknet_leaf_26_clk),
    .D(net1016),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7444_ (.CLK(clknet_leaf_40_clk),
    .D(net1236),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7445_ (.CLK(clknet_leaf_23_clk),
    .D(net1447),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7446_ (.CLK(clknet_leaf_22_clk),
    .D(net1058),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7447_ (.CLK(clknet_leaf_33_clk),
    .D(net1240),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7448_ (.CLK(clknet_leaf_25_clk),
    .D(net1170),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7449_ (.CLK(clknet_leaf_56_clk),
    .D(net1693),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7450_ (.CLK(clknet_leaf_28_clk),
    .D(net1232),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7451_ (.CLK(clknet_leaf_44_clk),
    .D(net1559),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7452_ (.CLK(clknet_leaf_21_clk),
    .D(net1318),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7453_ (.CLK(clknet_leaf_26_clk),
    .D(net1639),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7454_ (.CLK(clknet_leaf_49_clk),
    .D(net1358),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7455_ (.CLK(clknet_leaf_52_clk),
    .D(net968),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7456_ (.CLK(clknet_leaf_31_clk),
    .D(net1507),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7457_ (.CLK(clknet_leaf_50_clk),
    .D(net926),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7458_ (.CLK(clknet_leaf_54_clk),
    .D(net1362),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7459_ (.CLK(clknet_leaf_58_clk),
    .D(net1348),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7460_ (.CLK(clknet_leaf_47_clk),
    .D(net1056),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7461_ (.CLK(clknet_leaf_62_clk),
    .D(net1152),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7462_ (.CLK(clknet_leaf_30_clk),
    .D(net1040),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7463_ (.CLK(clknet_leaf_55_clk),
    .D(net1108),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7464_ (.CLK(clknet_leaf_60_clk),
    .D(net1354),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7465_ (.CLK(clknet_leaf_46_clk),
    .D(net1581),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7466_ (.CLK(clknet_leaf_53_clk),
    .D(net1024),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7467_ (.CLK(clknet_leaf_54_clk),
    .D(net1194),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7468_ (.CLK(clknet_leaf_29_clk),
    .D(net990),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7469_ (.CLK(clknet_leaf_43_clk),
    .D(net1180),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7470_ (.CLK(clknet_leaf_32_clk),
    .D(net904),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7471_ (.CLK(clknet_leaf_35_clk),
    .D(net1218),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7472_ (.CLK(clknet_leaf_40_clk),
    .D(net1202),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7473_ (.CLK(clknet_leaf_32_clk),
    .D(net813),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7474_ (.CLK(clknet_leaf_28_clk),
    .D(net1655),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7475_ (.CLK(clknet_leaf_24_clk),
    .D(net1034),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7476_ (.CLK(clknet_leaf_40_clk),
    .D(net1220),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7477_ (.CLK(clknet_leaf_48_clk),
    .D(net1555),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7478_ (.CLK(clknet_leaf_22_clk),
    .D(net1264),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7479_ (.CLK(clknet_leaf_35_clk),
    .D(net1366),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7480_ (.CLK(clknet_leaf_25_clk),
    .D(net1022),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7481_ (.CLK(clknet_leaf_56_clk),
    .D(net1621),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7482_ (.CLK(clknet_leaf_29_clk),
    .D(net935),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7483_ (.CLK(clknet_leaf_44_clk),
    .D(net1501),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7484_ (.CLK(clknet_leaf_23_clk),
    .D(net1425),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7485_ (.CLK(clknet_leaf_31_clk),
    .D(net1583),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7486_ (.CLK(clknet_leaf_49_clk),
    .D(net1288),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7487_ (.CLK(clknet_leaf_52_clk),
    .D(net998),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7488_ (.CLK(clknet_leaf_31_clk),
    .D(net1268),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7489_ (.CLK(clknet_leaf_49_clk),
    .D(net1441),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7490_ (.CLK(clknet_leaf_56_clk),
    .D(net1651),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7491_ (.CLK(clknet_leaf_58_clk),
    .D(net1038),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7492_ (.CLK(clknet_leaf_46_clk),
    .D(net1511),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7493_ (.CLK(clknet_leaf_60_clk),
    .D(net1681),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7494_ (.CLK(clknet_leaf_30_clk),
    .D(net1060),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7495_ (.CLK(clknet_leaf_56_clk),
    .D(net1687),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7496_ (.CLK(clknet_leaf_60_clk),
    .D(net1615),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7497_ (.CLK(clknet_leaf_42_clk),
    .D(net1304),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7498_ (.CLK(clknet_leaf_56_clk),
    .D(net1370),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7499_ (.CLK(clknet_leaf_54_clk),
    .D(net1827),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7500_ (.CLK(clknet_leaf_30_clk),
    .D(net939),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7501_ (.CLK(clknet_leaf_43_clk),
    .D(net1286),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7502_ (.CLK(net480),
    .D(_0000_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7503_ (.CLK(net481),
    .D(_0011_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7504_ (.CLK(net482),
    .D(_0022_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7505_ (.CLK(net483),
    .D(_0025_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7506_ (.CLK(net484),
    .D(_0026_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7507_ (.CLK(net485),
    .D(_0027_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7508_ (.CLK(net486),
    .D(_0028_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7509_ (.CLK(net487),
    .D(_0029_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7510_ (.CLK(net488),
    .D(_0030_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7511_ (.CLK(net489),
    .D(_0031_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7512_ (.CLK(net490),
    .D(_0001_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7513_ (.CLK(net491),
    .D(_0002_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7514_ (.CLK(net492),
    .D(_0003_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7515_ (.CLK(net493),
    .D(_0004_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7516_ (.CLK(net494),
    .D(_0005_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7517_ (.CLK(net495),
    .D(_0006_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7518_ (.CLK(net496),
    .D(_0007_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7519_ (.CLK(net497),
    .D(_0008_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7520_ (.CLK(net498),
    .D(_0009_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7521_ (.CLK(net499),
    .D(_0010_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7522_ (.CLK(net500),
    .D(_0012_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7523_ (.CLK(net501),
    .D(_0013_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7524_ (.CLK(net502),
    .D(_0014_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7525_ (.CLK(net503),
    .D(_0015_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7526_ (.CLK(net504),
    .D(_0016_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7527_ (.CLK(net505),
    .D(_0017_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7528_ (.CLK(net506),
    .D(_0018_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7529_ (.CLK(net507),
    .D(_0019_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7530_ (.CLK(net508),
    .D(_0020_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7531_ (.CLK(net509),
    .D(_0021_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7532_ (.CLK(net510),
    .D(_0023_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7533_ (.CLK(net511),
    .D(_0024_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7534_ (.CLK(clknet_leaf_38_clk),
    .D(net1605),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7535_ (.CLK(clknet_leaf_38_clk),
    .D(net1661),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7536_ (.CLK(clknet_leaf_39_clk),
    .D(net802),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7537_ (.CLK(clknet_leaf_38_clk),
    .D(net914),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7538_ (.CLK(clknet_leaf_27_clk),
    .D(net1004),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7539_ (.CLK(clknet_leaf_25_clk),
    .D(net1503),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7540_ (.CLK(clknet_leaf_46_clk),
    .D(net1479),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7541_ (.CLK(clknet_leaf_23_clk),
    .D(net1262),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7542_ (.CLK(clknet_leaf_22_clk),
    .D(net1112),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7543_ (.CLK(clknet_leaf_33_clk),
    .D(net1132),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7544_ (.CLK(clknet_leaf_25_clk),
    .D(net1346),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7545_ (.CLK(clknet_leaf_57_clk),
    .D(net1176),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7546_ (.CLK(clknet_leaf_27_clk),
    .D(net1014),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7547_ (.CLK(clknet_leaf_44_clk),
    .D(net1619),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7548_ (.CLK(clknet_leaf_21_clk),
    .D(net1328),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7549_ (.CLK(clknet_leaf_26_clk),
    .D(net1160),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7550_ (.CLK(clknet_leaf_49_clk),
    .D(net1000),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7551_ (.CLK(clknet_leaf_52_clk),
    .D(net1106),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7552_ (.CLK(clknet_leaf_31_clk),
    .D(net1400),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7553_ (.CLK(clknet_leaf_21_clk),
    .D(net1284),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7554_ (.CLK(clknet_leaf_54_clk),
    .D(net1467),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7555_ (.CLK(clknet_leaf_57_clk),
    .D(net1368),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7556_ (.CLK(clknet_leaf_47_clk),
    .D(net1044),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7557_ (.CLK(clknet_leaf_56_clk),
    .D(net1412),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7558_ (.CLK(clknet_leaf_31_clk),
    .D(net1320),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7559_ (.CLK(clknet_leaf_56_clk),
    .D(net1669),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7560_ (.CLK(clknet_leaf_58_clk),
    .D(net1527),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7561_ (.CLK(clknet_leaf_46_clk),
    .D(net1280),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7562_ (.CLK(clknet_leaf_53_clk),
    .D(net953),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7563_ (.CLK(clknet_leaf_54_clk),
    .D(net1178),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7564_ (.CLK(clknet_leaf_31_clk),
    .D(net1374),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7565_ (.CLK(clknet_leaf_57_clk),
    .D(net1292),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7566_ (.CLK(clknet_leaf_38_clk),
    .D(net853),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7567_ (.CLK(clknet_leaf_38_clk),
    .D(net1775),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7568_ (.CLK(clknet_leaf_38_clk),
    .D(net1098),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7569_ (.CLK(clknet_leaf_38_clk),
    .D(net955),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7570_ (.CLK(clknet_leaf_27_clk),
    .D(net1156),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7571_ (.CLK(clknet_leaf_25_clk),
    .D(net1585),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7572_ (.CLK(clknet_leaf_39_clk),
    .D(net1324),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7573_ (.CLK(clknet_leaf_23_clk),
    .D(net1258),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7574_ (.CLK(clknet_leaf_22_clk),
    .D(net951),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7575_ (.CLK(clknet_leaf_33_clk),
    .D(net1338),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7576_ (.CLK(clknet_leaf_25_clk),
    .D(net1248),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7577_ (.CLK(clknet_leaf_57_clk),
    .D(net1196),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7578_ (.CLK(clknet_leaf_27_clk),
    .D(net924),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7579_ (.CLK(clknet_leaf_44_clk),
    .D(net1519),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7580_ (.CLK(clknet_leaf_21_clk),
    .D(net1356),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7581_ (.CLK(clknet_leaf_26_clk),
    .D(net1050),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7582_ (.CLK(clknet_leaf_49_clk),
    .D(net1224),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7583_ (.CLK(clknet_leaf_52_clk),
    .D(net1002),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7584_ (.CLK(clknet_leaf_31_clk),
    .D(net1410),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7585_ (.CLK(clknet_leaf_21_clk),
    .D(net1475),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7586_ (.CLK(clknet_leaf_56_clk),
    .D(net1408),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7587_ (.CLK(clknet_leaf_57_clk),
    .D(net1064),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7588_ (.CLK(clknet_leaf_48_clk),
    .D(net1495),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7589_ (.CLK(clknet_leaf_56_clk),
    .D(net1308),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7590_ (.CLK(clknet_leaf_31_clk),
    .D(net1419),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7591_ (.CLK(clknet_leaf_56_clk),
    .D(net1300),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7592_ (.CLK(clknet_leaf_56_clk),
    .D(net1392),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7593_ (.CLK(clknet_leaf_46_clk),
    .D(net1719),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7594_ (.CLK(clknet_leaf_57_clk),
    .D(net1254),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7595_ (.CLK(clknet_leaf_54_clk),
    .D(net1449),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7596_ (.CLK(clknet_leaf_31_clk),
    .D(net1675),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7597_ (.CLK(clknet_leaf_57_clk),
    .D(net1084),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7598_ (.CLK(clknet_leaf_38_clk),
    .D(net1729),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7599_ (.CLK(clknet_leaf_33_clk),
    .D(net1671),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7600_ (.CLK(clknet_leaf_39_clk),
    .D(net791),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7601_ (.CLK(clknet_leaf_39_clk),
    .D(net1934),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7602_ (.CLK(clknet_leaf_29_clk),
    .D(net1070),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7603_ (.CLK(clknet_leaf_25_clk),
    .D(net1396),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7604_ (.CLK(clknet_leaf_40_clk),
    .D(net1543),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7605_ (.CLK(clknet_leaf_23_clk),
    .D(net1551),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7606_ (.CLK(clknet_leaf_22_clk),
    .D(net1230),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7607_ (.CLK(clknet_leaf_33_clk),
    .D(net1350),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7608_ (.CLK(clknet_leaf_24_clk),
    .D(net1234),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7609_ (.CLK(clknet_leaf_57_clk),
    .D(net1635),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7610_ (.CLK(clknet_leaf_31_clk),
    .D(net1433),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7611_ (.CLK(clknet_leaf_43_clk),
    .D(net1653),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7612_ (.CLK(clknet_leaf_23_clk),
    .D(net1805),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7613_ (.CLK(clknet_leaf_27_clk),
    .D(net1571),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7614_ (.CLK(clknet_leaf_45_clk),
    .D(net1256),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7615_ (.CLK(clknet_leaf_54_clk),
    .D(net1695),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7616_ (.CLK(clknet_leaf_31_clk),
    .D(net1691),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7617_ (.CLK(clknet_leaf_50_clk),
    .D(net1172),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7618_ (.CLK(clknet_leaf_56_clk),
    .D(net1469),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7619_ (.CLK(clknet_leaf_58_clk),
    .D(net1633),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7620_ (.CLK(clknet_leaf_46_clk),
    .D(net1535),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7621_ (.CLK(clknet_leaf_60_clk),
    .D(net1625),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7622_ (.CLK(clknet_leaf_33_clk),
    .D(net1326),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7623_ (.CLK(clknet_leaf_58_clk),
    .D(net1579),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7624_ (.CLK(clknet_leaf_60_clk),
    .D(net1641),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7625_ (.CLK(clknet_leaf_44_clk),
    .D(net1250),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7626_ (.CLK(clknet_leaf_56_clk),
    .D(net1645),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7627_ (.CLK(clknet_leaf_56_clk),
    .D(net1815),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7628_ (.CLK(clknet_leaf_31_clk),
    .D(net1611),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7629_ (.CLK(clknet_leaf_58_clk),
    .D(net1330),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7630_ (.CLK(clknet_leaf_2_clk),
    .D(_0507_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_src_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7631_ (.CLK(clknet_leaf_78_clk),
    .D(_0508_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7632_ (.CLK(clknet_leaf_2_clk),
    .D(_0509_),
    .Q(\U_DATAPATH.U_EX_MEM.i_mem_write_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7633_ (.CLK(clknet_leaf_2_clk),
    .D(_0510_),
    .Q(\U_DATAPATH.U_EX_MEM.i_result_src_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7634_ (.CLK(clknet_leaf_17_clk),
    .D(_0511_),
    .Q(\U_DATAPATH.U_EX_MEM.i_reg_write_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7635_ (.CLK(clknet_leaf_73_clk),
    .D(net1118),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7636_ (.CLK(clknet_leaf_16_clk),
    .D(net895),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7637_ (.CLK(clknet_leaf_16_clk),
    .D(net839),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7638_ (.CLK(clknet_leaf_7_clk),
    .D(net887),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7639_ (.CLK(clknet_leaf_17_clk),
    .D(net883),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7640_ (.CLK(clknet_leaf_15_clk),
    .D(net931),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7641_ (.CLK(clknet_leaf_15_clk),
    .D(net763),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7642_ (.CLK(clknet_leaf_15_clk),
    .D(net920),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7643_ (.CLK(clknet_leaf_6_clk),
    .D(net902),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7644_ (.CLK(clknet_leaf_6_clk),
    .D(net833),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7645_ (.CLK(clknet_leaf_15_clk),
    .D(net835),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7646_ (.CLK(clknet_leaf_19_clk),
    .D(net808),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7647_ (.CLK(clknet_leaf_6_clk),
    .D(net1042),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7648_ (.CLK(clknet_leaf_6_clk),
    .D(net857),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7649_ (.CLK(clknet_leaf_48_clk),
    .D(net1030),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7650_ (.CLK(clknet_leaf_21_clk),
    .D(net609),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7651_ (.CLK(clknet_leaf_47_clk),
    .D(net1032),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7652_ (.CLK(clknet_leaf_52_clk),
    .D(net800),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7653_ (.CLK(clknet_leaf_75_clk),
    .D(net1126),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7654_ (.CLK(clknet_leaf_64_clk),
    .D(net872),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7655_ (.CLK(clknet_leaf_69_clk),
    .D(net949),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7656_ (.CLK(clknet_leaf_64_clk),
    .D(net916),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7657_ (.CLK(clknet_leaf_69_clk),
    .D(net821),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7658_ (.CLK(clknet_leaf_66_clk),
    .D(net775),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7659_ (.CLK(clknet_leaf_64_clk),
    .D(net765),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7660_ (.CLK(clknet_leaf_66_clk),
    .D(net804),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7661_ (.CLK(clknet_leaf_72_clk),
    .D(net984),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7662_ (.CLK(clknet_leaf_72_clk),
    .D(net659),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7663_ (.CLK(clknet_leaf_72_clk),
    .D(net1282),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7664_ (.CLK(clknet_leaf_67_clk),
    .D(net773),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7665_ (.CLK(clknet_leaf_72_clk),
    .D(net555),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7666_ (.CLK(clknet_leaf_18_clk),
    .D(net1136),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7667_ (.CLK(clknet_leaf_18_clk),
    .D(net970),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7668_ (.CLK(clknet_leaf_17_clk),
    .D(net726),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7669_ (.CLK(clknet_leaf_19_clk),
    .D(net843),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7670_ (.CLK(clknet_leaf_7_clk),
    .D(net841),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7671_ (.CLK(clknet_leaf_16_clk),
    .D(net742),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7672_ (.CLK(clknet_leaf_14_clk),
    .D(net789),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7673_ (.CLK(clknet_leaf_4_clk),
    .D(net553),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7674_ (.CLK(clknet_leaf_5_clk),
    .D(net823),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7675_ (.CLK(clknet_leaf_13_clk),
    .D(net581),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7676_ (.CLK(clknet_leaf_49_clk),
    .D(net879),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7677_ (.CLK(clknet_leaf_19_clk),
    .D(net885),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7678_ (.CLK(clknet_leaf_13_clk),
    .D(net793),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7679_ (.CLK(clknet_leaf_50_clk),
    .D(net549),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7680_ (.CLK(clknet_leaf_48_clk),
    .D(net1228),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7681_ (.CLK(clknet_leaf_14_clk),
    .D(net1078),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7682_ (.CLK(clknet_leaf_57_clk),
    .D(net1096),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7683_ (.CLK(clknet_leaf_71_clk),
    .D(net849),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7684_ (.CLK(clknet_leaf_63_clk),
    .D(net1062),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7685_ (.CLK(clknet_leaf_63_clk),
    .D(net1018),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7686_ (.CLK(clknet_leaf_67_clk),
    .D(net910),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7687_ (.CLK(clknet_leaf_64_clk),
    .D(net961),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7688_ (.CLK(clknet_leaf_67_clk),
    .D(net957),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7689_ (.CLK(clknet_leaf_68_clk),
    .D(net1086),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7690_ (.CLK(clknet_leaf_68_clk),
    .D(net649),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7691_ (.CLK(clknet_leaf_71_clk),
    .D(net876),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7692_ (.CLK(clknet_leaf_72_clk),
    .D(net1066),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7693_ (.CLK(clknet_leaf_70_clk),
    .D(net815),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7694_ (.CLK(clknet_leaf_67_clk),
    .D(net864),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7695_ (.CLK(clknet_leaf_32_clk),
    .D(_0572_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7696_ (.CLK(clknet_leaf_32_clk),
    .D(_0573_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7697_ (.CLK(clknet_leaf_24_clk),
    .D(_0574_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7698_ (.CLK(clknet_leaf_32_clk),
    .D(_0575_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7699_ (.CLK(clknet_leaf_39_clk),
    .D(_0576_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7700_ (.CLK(clknet_leaf_47_clk),
    .D(_0577_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7701_ (.CLK(clknet_leaf_46_clk),
    .D(_0578_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7702_ (.CLK(clknet_leaf_47_clk),
    .D(_0579_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7703_ (.CLK(clknet_leaf_39_clk),
    .D(_0580_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7704_ (.CLK(clknet_leaf_33_clk),
    .D(_0581_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7705_ (.CLK(clknet_leaf_45_clk),
    .D(_0582_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7706_ (.CLK(clknet_leaf_33_clk),
    .D(_0583_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7707_ (.CLK(clknet_leaf_13_clk),
    .D(_0584_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7708_ (.CLK(clknet_leaf_22_clk),
    .D(_0585_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7709_ (.CLK(clknet_leaf_46_clk),
    .D(_0586_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7710_ (.CLK(clknet_leaf_48_clk),
    .D(_0587_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7711_ (.CLK(clknet_leaf_18_clk),
    .D(_0588_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7712_ (.CLK(clknet_leaf_13_clk),
    .D(_0589_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7713_ (.CLK(clknet_leaf_21_clk),
    .D(_0590_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7714_ (.CLK(clknet_leaf_56_clk),
    .D(_0591_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7715_ (.CLK(clknet_leaf_13_clk),
    .D(_0592_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7716_ (.CLK(clknet_leaf_44_clk),
    .D(_0593_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7717_ (.CLK(clknet_leaf_20_clk),
    .D(_0594_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7718_ (.CLK(clknet_leaf_13_clk),
    .D(_0595_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7719_ (.CLK(clknet_leaf_45_clk),
    .D(_0596_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7720_ (.CLK(clknet_leaf_76_clk),
    .D(_0597_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7721_ (.CLK(clknet_leaf_24_clk),
    .D(_0598_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7722_ (.CLK(clknet_leaf_51_clk),
    .D(_0599_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7723_ (.CLK(clknet_leaf_55_clk),
    .D(_0600_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7724_ (.CLK(clknet_leaf_61_clk),
    .D(_0601_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7725_ (.CLK(clknet_leaf_48_clk),
    .D(_0602_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7726_ (.CLK(clknet_leaf_64_clk),
    .D(_0603_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7727_ (.CLK(clknet_leaf_31_clk),
    .D(_0604_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7728_ (.CLK(clknet_leaf_62_clk),
    .D(_0605_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7729_ (.CLK(clknet_leaf_65_clk),
    .D(_0606_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7730_ (.CLK(clknet_leaf_44_clk),
    .D(_0607_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7731_ (.CLK(clknet_leaf_75_clk),
    .D(_0608_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7732_ (.CLK(clknet_leaf_75_clk),
    .D(_0609_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7733_ (.CLK(clknet_leaf_31_clk),
    .D(_0610_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7734_ (.CLK(clknet_leaf_61_clk),
    .D(_0611_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7735_ (.CLK(clknet_leaf_42_clk),
    .D(_0612_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7736_ (.CLK(clknet_leaf_33_clk),
    .D(_0613_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7737_ (.CLK(clknet_leaf_46_clk),
    .D(_0614_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7738_ (.CLK(clknet_leaf_32_clk),
    .D(_0615_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7739_ (.CLK(clknet_leaf_13_clk),
    .D(_0616_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7740_ (.CLK(clknet_leaf_13_clk),
    .D(_0617_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7741_ (.CLK(clknet_leaf_46_clk),
    .D(_0618_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7742_ (.CLK(clknet_leaf_21_clk),
    .D(_0619_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7743_ (.CLK(clknet_leaf_18_clk),
    .D(_0620_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7744_ (.CLK(clknet_leaf_12_clk),
    .D(_0621_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7745_ (.CLK(clknet_leaf_14_clk),
    .D(_0622_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7746_ (.CLK(clknet_leaf_77_clk),
    .D(_0623_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7747_ (.CLK(clknet_leaf_13_clk),
    .D(_0624_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7748_ (.CLK(clknet_leaf_44_clk),
    .D(_0625_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7749_ (.CLK(clknet_leaf_20_clk),
    .D(_0626_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7750_ (.CLK(clknet_leaf_13_clk),
    .D(_0627_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7751_ (.CLK(clknet_leaf_49_clk),
    .D(_0628_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7752_ (.CLK(clknet_leaf_54_clk),
    .D(_0629_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7753_ (.CLK(clknet_leaf_24_clk),
    .D(_0630_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7754_ (.CLK(clknet_leaf_51_clk),
    .D(_0631_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7755_ (.CLK(clknet_leaf_55_clk),
    .D(_0632_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7756_ (.CLK(clknet_leaf_65_clk),
    .D(_0633_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7757_ (.CLK(clknet_leaf_63_clk),
    .D(_0634_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7758_ (.CLK(clknet_leaf_65_clk),
    .D(_0635_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[23] ));
 sky130_fd_sc_hd__dfxtp_4 _7759_ (.CLK(clknet_leaf_32_clk),
    .D(_0636_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7760_ (.CLK(clknet_leaf_64_clk),
    .D(_0637_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7761_ (.CLK(clknet_leaf_64_clk),
    .D(_0638_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7762_ (.CLK(clknet_leaf_65_clk),
    .D(_0639_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7763_ (.CLK(clknet_leaf_69_clk),
    .D(_0640_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7764_ (.CLK(clknet_leaf_69_clk),
    .D(_0641_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[29] ));
 sky130_fd_sc_hd__dfxtp_4 _7765_ (.CLK(clknet_leaf_31_clk),
    .D(_0642_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7766_ (.CLK(clknet_leaf_65_clk),
    .D(_0643_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7767_ (.CLK(clknet_leaf_18_clk),
    .D(_0644_),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7768_ (.CLK(clknet_leaf_18_clk),
    .D(_0645_),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7769_ (.CLK(clknet_leaf_22_clk),
    .D(_0646_),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7770_ (.CLK(clknet_leaf_22_clk),
    .D(net2108),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ));
 sky130_fd_sc_hd__dfxtp_2 _7771_ (.CLK(clknet_leaf_2_clk),
    .D(_0648_),
    .Q(\U_DATAPATH.U_ID_EX.o_addr_src_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7772_ (.CLK(clknet_leaf_1_clk),
    .D(_0649_),
    .Q(\U_CONTROL_UNIT.i_branch_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7773_ (.CLK(clknet_leaf_1_clk),
    .D(_0650_),
    .Q(\U_CONTROL_UNIT.i_jump_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7774_ (.CLK(clknet_leaf_50_clk),
    .D(net1880),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7775_ (.CLK(clknet_leaf_51_clk),
    .D(net2139),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7776_ (.CLK(clknet_leaf_72_clk),
    .D(_0653_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7777_ (.CLK(clknet_leaf_17_clk),
    .D(_0654_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7778_ (.CLK(clknet_leaf_17_clk),
    .D(_0655_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7779_ (.CLK(clknet_leaf_17_clk),
    .D(_0656_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7780_ (.CLK(clknet_leaf_18_clk),
    .D(_0657_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7781_ (.CLK(clknet_leaf_14_clk),
    .D(_0658_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7782_ (.CLK(clknet_leaf_15_clk),
    .D(_0659_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7783_ (.CLK(clknet_leaf_14_clk),
    .D(_0660_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7784_ (.CLK(clknet_leaf_7_clk),
    .D(_0661_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7785_ (.CLK(clknet_leaf_4_clk),
    .D(_0662_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7786_ (.CLK(clknet_leaf_15_clk),
    .D(_0663_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7787_ (.CLK(clknet_leaf_4_clk),
    .D(_0664_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7788_ (.CLK(clknet_leaf_5_clk),
    .D(_0665_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7789_ (.CLK(clknet_leaf_4_clk),
    .D(_0666_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7790_ (.CLK(clknet_leaf_48_clk),
    .D(_0667_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7791_ (.CLK(clknet_leaf_50_clk),
    .D(_0668_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7792_ (.CLK(clknet_leaf_24_clk),
    .D(_0669_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7793_ (.CLK(clknet_leaf_53_clk),
    .D(_0670_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7794_ (.CLK(clknet_leaf_55_clk),
    .D(_0671_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7795_ (.CLK(clknet_leaf_64_clk),
    .D(_0672_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7796_ (.CLK(clknet_leaf_75_clk),
    .D(_0673_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7797_ (.CLK(clknet_leaf_64_clk),
    .D(_0674_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7798_ (.CLK(clknet_leaf_68_clk),
    .D(_0675_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7799_ (.CLK(clknet_leaf_68_clk),
    .D(_0676_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7800_ (.CLK(clknet_leaf_64_clk),
    .D(_0677_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7801_ (.CLK(clknet_leaf_66_clk),
    .D(_0678_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7802_ (.CLK(clknet_leaf_70_clk),
    .D(_0679_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7803_ (.CLK(clknet_leaf_70_clk),
    .D(_0680_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7804_ (.CLK(clknet_leaf_70_clk),
    .D(_0681_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7805_ (.CLK(clknet_leaf_67_clk),
    .D(_0682_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7806_ (.CLK(clknet_leaf_47_clk),
    .D(net2010),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7807_ (.CLK(clknet_leaf_47_clk),
    .D(net1869),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7808_ (.CLK(clknet_leaf_47_clk),
    .D(net661),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7809_ (.CLK(clknet_leaf_47_clk),
    .D(net744),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7810_ (.CLK(clknet_leaf_72_clk),
    .D(net547),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7811_ (.CLK(clknet_leaf_16_clk),
    .D(net667),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7812_ (.CLK(clknet_leaf_17_clk),
    .D(net583),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7813_ (.CLK(clknet_leaf_16_clk),
    .D(net589),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7814_ (.CLK(clknet_leaf_19_clk),
    .D(net601),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7815_ (.CLK(clknet_leaf_14_clk),
    .D(net603),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7816_ (.CLK(clknet_leaf_15_clk),
    .D(net714),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7817_ (.CLK(clknet_leaf_15_clk),
    .D(net708),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7818_ (.CLK(clknet_leaf_6_clk),
    .D(net680),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7819_ (.CLK(clknet_leaf_2_clk),
    .D(net781),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7820_ (.CLK(clknet_leaf_15_clk),
    .D(net732),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7821_ (.CLK(clknet_leaf_4_clk),
    .D(net577),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7822_ (.CLK(clknet_leaf_6_clk),
    .D(net678),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7823_ (.CLK(clknet_leaf_5_clk),
    .D(net615),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7824_ (.CLK(clknet_leaf_48_clk),
    .D(net696),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7825_ (.CLK(clknet_leaf_21_clk),
    .D(net730),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7826_ (.CLK(clknet_leaf_47_clk),
    .D(net698),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7827_ (.CLK(clknet_leaf_53_clk),
    .D(net567),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7828_ (.CLK(clknet_leaf_63_clk),
    .D(net557),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7829_ (.CLK(clknet_leaf_64_clk),
    .D(net716),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7830_ (.CLK(clknet_leaf_69_clk),
    .D(net718),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7831_ (.CLK(clknet_leaf_64_clk),
    .D(net753),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7832_ (.CLK(clknet_leaf_69_clk),
    .D(net692),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7833_ (.CLK(clknet_leaf_66_clk),
    .D(net651),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7834_ (.CLK(clknet_leaf_65_clk),
    .D(net637),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7835_ (.CLK(clknet_leaf_66_clk),
    .D(net657),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7836_ (.CLK(clknet_leaf_72_clk),
    .D(net738),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7837_ (.CLK(clknet_leaf_72_clk),
    .D(net755),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7838_ (.CLK(clknet_leaf_72_clk),
    .D(net757),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7839_ (.CLK(clknet_leaf_67_clk),
    .D(net736),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[31] ));
 sky130_fd_sc_hd__dfxtp_2 _7840_ (.CLK(clknet_leaf_4_clk),
    .D(_0717_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_4 _7841_ (.CLK(clknet_leaf_77_clk),
    .D(_0718_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_4 _7842_ (.CLK(clknet_leaf_76_clk),
    .D(_0719_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_4 _7843_ (.CLK(clknet_leaf_78_clk),
    .D(_0720_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_2 _7844_ (.CLK(clknet_leaf_77_clk),
    .D(_0721_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_2 _7845_ (.CLK(clknet_leaf_18_clk),
    .D(_0722_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_4 _7846_ (.CLK(clknet_leaf_3_clk),
    .D(_0723_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_4 _7847_ (.CLK(clknet_leaf_80_clk),
    .D(_0724_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_4 _7848_ (.CLK(clknet_leaf_78_clk),
    .D(_0725_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_4 _7849_ (.CLK(clknet_leaf_78_clk),
    .D(net2338),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_2 _7850_ (.CLK(clknet_leaf_3_clk),
    .D(_0727_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_4 _7851_ (.CLK(clknet_leaf_80_clk),
    .D(_0728_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_4 _7852_ (.CLK(clknet_leaf_3_clk),
    .D(net2290),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_4 _7853_ (.CLK(clknet_leaf_52_clk),
    .D(net2315),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_4 _7854_ (.CLK(clknet_leaf_19_clk),
    .D(net2322),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_2 _7855_ (.CLK(clknet_leaf_18_clk),
    .D(_0732_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_4 _7856_ (.CLK(clknet_leaf_52_clk),
    .D(net2304),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_2 _7857_ (.CLK(clknet_leaf_76_clk),
    .D(net2306),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_4 _7858_ (.CLK(clknet_leaf_20_clk),
    .D(_0735_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_4 _7859_ (.CLK(clknet_leaf_51_clk),
    .D(_0736_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_2 _7860_ (.CLK(clknet_leaf_75_clk),
    .D(_0737_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_2 _7861_ (.CLK(clknet_leaf_75_clk),
    .D(net2311),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_4 _7862_ (.CLK(clknet_leaf_75_clk),
    .D(net2296),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_2 _7863_ (.CLK(clknet_leaf_74_clk),
    .D(net2308),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_4 _7864_ (.CLK(clknet_leaf_74_clk),
    .D(_0741_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_4 _7865_ (.CLK(clknet_leaf_73_clk),
    .D(net2285),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_2 _7866_ (.CLK(clknet_leaf_68_clk),
    .D(_0743_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_2 _7867_ (.CLK(clknet_leaf_69_clk),
    .D(net2332),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_4 _7868_ (.CLK(clknet_leaf_81_clk),
    .D(net2272),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_4 _7869_ (.CLK(clknet_leaf_72_clk),
    .D(net2262),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_4 _7870_ (.CLK(clknet_leaf_78_clk),
    .D(_0747_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_4 _7871_ (.CLK(clknet_leaf_70_clk),
    .D(_0748_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _7872_ (.CLK(clknet_leaf_3_clk),
    .D(_0749_),
    .Q(\U_DATAPATH.U_EX_MEM.o_result_src_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7873_ (.CLK(clknet_leaf_4_clk),
    .D(net611),
    .Q(\U_DATAPATH.U_EX_MEM.o_result_src_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7874_ (.CLK(clknet_leaf_47_clk),
    .D(net740),
    .Q(\U_DATAPATH.U_EX_MEM.o_reg_write_M ));
 sky130_fd_sc_hd__dfxtp_2 _7875_ (.CLK(clknet_leaf_60_clk),
    .D(_0752_),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_1 _7876_ (.CLK(clknet_leaf_83_clk),
    .D(_0753_),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_1 _7877_ (.CLK(clknet_leaf_84_clk),
    .D(_0754_),
    .Q(net152));
 sky130_fd_sc_hd__dfxtp_1 _7878_ (.CLK(clknet_leaf_34_clk),
    .D(_0755_),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_1 _7879_ (.CLK(clknet_leaf_28_clk),
    .D(_0756_),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_2 _7880_ (.CLK(clknet_leaf_13_clk),
    .D(_0757_),
    .Q(net157));
 sky130_fd_sc_hd__dfxtp_2 _7881_ (.CLK(clknet_leaf_13_clk),
    .D(_0758_),
    .Q(net158));
 sky130_fd_sc_hd__dfxtp_2 _7882_ (.CLK(clknet_leaf_59_clk),
    .D(_0759_),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_1 _7883_ (.CLK(clknet_leaf_79_clk),
    .D(_0760_),
    .Q(net160));
 sky130_fd_sc_hd__dfxtp_1 _7884_ (.CLK(clknet_3_4_0_clk),
    .D(_0761_),
    .Q(net161));
 sky130_fd_sc_hd__dfxtp_2 _7885_ (.CLK(clknet_leaf_41_clk),
    .D(_0762_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_2 _7886_ (.CLK(clknet_leaf_79_clk),
    .D(_0763_),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_1 _7887_ (.CLK(clknet_leaf_6_clk),
    .D(_0764_),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_1 _7888_ (.CLK(clknet_leaf_66_clk),
    .D(_0765_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_2 _7889_ (.CLK(clknet_leaf_78_clk),
    .D(_0766_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_1 _7890_ (.CLK(clknet_leaf_81_clk),
    .D(_0767_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_1 _7891_ (.CLK(clknet_leaf_9_clk),
    .D(_0768_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_2 _7892_ (.CLK(clknet_leaf_0_clk),
    .D(net2254),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_1 _7893_ (.CLK(clknet_leaf_12_clk),
    .D(_0770_),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_1 _7894_ (.CLK(clknet_leaf_9_clk),
    .D(_0771_),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_2 _7895_ (.CLK(clknet_leaf_84_clk),
    .D(_0772_),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_2 _7896_ (.CLK(clknet_leaf_72_clk),
    .D(_0773_),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_1 _7897_ (.CLK(clknet_leaf_12_clk),
    .D(_0774_),
    .Q(net144));
 sky130_fd_sc_hd__dfxtp_1 _7898_ (.CLK(clknet_leaf_71_clk),
    .D(_0775_),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_1 _7899_ (.CLK(clknet_leaf_35_clk),
    .D(_0776_),
    .Q(net146));
 sky130_fd_sc_hd__dfxtp_1 _7900_ (.CLK(clknet_leaf_61_clk),
    .D(_0777_),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_2 _7901_ (.CLK(clknet_leaf_72_clk),
    .D(_0778_),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_1 _7902_ (.CLK(clknet_leaf_41_clk),
    .D(_0779_),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_1 _7903_ (.CLK(clknet_leaf_82_clk),
    .D(_0780_),
    .Q(net150));
 sky130_fd_sc_hd__dfxtp_1 _7904_ (.CLK(clknet_leaf_73_clk),
    .D(_0781_),
    .Q(net151));
 sky130_fd_sc_hd__dfxtp_1 _7905_ (.CLK(clknet_leaf_41_clk),
    .D(_0782_),
    .Q(net153));
 sky130_fd_sc_hd__dfxtp_1 _7906_ (.CLK(clknet_leaf_66_clk),
    .D(_0783_),
    .Q(net154));
 sky130_fd_sc_hd__dfxtp_2 _7907_ (.CLK(clknet_leaf_0_clk),
    .D(_0784_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_1 _7908_ (.CLK(clknet_leaf_28_clk),
    .D(net597),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _7909_ (.CLK(clknet_leaf_28_clk),
    .D(net749),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_1 _7910_ (.CLK(clknet_leaf_83_clk),
    .D(_0787_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _7911_ (.CLK(clknet_leaf_47_clk),
    .D(_0788_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ));
 sky130_fd_sc_hd__dfxtp_2 _7912_ (.CLK(clknet_leaf_39_clk),
    .D(net2063),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7913_ (.CLK(clknet_leaf_47_clk),
    .D(net2039),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ));
 sky130_fd_sc_hd__dfxtp_4 _7914_ (.CLK(clknet_leaf_32_clk),
    .D(net1983),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ));
 sky130_fd_sc_hd__dfxtp_4 _7915_ (.CLK(clknet_leaf_32_clk),
    .D(net1986),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7916_ (.CLK(clknet_leaf_72_clk),
    .D(net771),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7917_ (.CLK(clknet_leaf_17_clk),
    .D(net587),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7918_ (.CLK(clknet_leaf_14_clk),
    .D(net627),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7919_ (.CLK(clknet_leaf_17_clk),
    .D(net585),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7920_ (.CLK(clknet_leaf_19_clk),
    .D(net690),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7921_ (.CLK(clknet_leaf_14_clk),
    .D(net734),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7922_ (.CLK(clknet_leaf_15_clk),
    .D(net710),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7923_ (.CLK(clknet_leaf_14_clk),
    .D(net599),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7924_ (.CLK(clknet_leaf_5_clk),
    .D(net625),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7925_ (.CLK(clknet_leaf_3_clk),
    .D(net653),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7926_ (.CLK(clknet_leaf_15_clk),
    .D(net751),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7927_ (.CLK(clknet_leaf_20_clk),
    .D(net605),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7928_ (.CLK(clknet_leaf_5_clk),
    .D(net619),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7929_ (.CLK(clknet_leaf_4_clk),
    .D(net575),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7930_ (.CLK(clknet_leaf_45_clk),
    .D(net663),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7931_ (.CLK(clknet_leaf_21_clk),
    .D(net728),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7932_ (.CLK(clknet_leaf_24_clk),
    .D(net565),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7933_ (.CLK(clknet_leaf_53_clk),
    .D(net706),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7934_ (.CLK(clknet_leaf_63_clk),
    .D(net655),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7935_ (.CLK(clknet_leaf_65_clk),
    .D(net629),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7936_ (.CLK(clknet_leaf_69_clk),
    .D(net682),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7937_ (.CLK(clknet_leaf_64_clk),
    .D(net702),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7938_ (.CLK(clknet_leaf_69_clk),
    .D(net724),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7939_ (.CLK(clknet_leaf_66_clk),
    .D(net700),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7940_ (.CLK(clknet_leaf_65_clk),
    .D(net684),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7941_ (.CLK(clknet_leaf_65_clk),
    .D(net593),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7942_ (.CLK(clknet_leaf_72_clk),
    .D(net769),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7943_ (.CLK(clknet_leaf_70_clk),
    .D(net1477),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[29] ));
 sky130_fd_sc_hd__dfxtp_2 _7944_ (.CLK(clknet_leaf_72_clk),
    .D(net767),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7945_ (.CLK(clknet_leaf_66_clk),
    .D(net595),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7946_ (.CLK(clknet_leaf_49_clk),
    .D(net569),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7947_ (.CLK(clknet_leaf_52_clk),
    .D(net551),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7948_ (.CLK(clknet_leaf_72_clk),
    .D(net747),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7949_ (.CLK(clknet_leaf_17_clk),
    .D(net704),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7950_ (.CLK(clknet_leaf_14_clk),
    .D(net623),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7951_ (.CLK(clknet_leaf_17_clk),
    .D(net676),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7952_ (.CLK(clknet_leaf_19_clk),
    .D(net617),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7953_ (.CLK(clknet_leaf_14_clk),
    .D(net722),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7954_ (.CLK(clknet_leaf_14_clk),
    .D(net613),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7955_ (.CLK(clknet_leaf_14_clk),
    .D(net674),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7956_ (.CLK(clknet_leaf_5_clk),
    .D(net573),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7957_ (.CLK(clknet_leaf_4_clk),
    .D(net688),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7958_ (.CLK(clknet_leaf_14_clk),
    .D(net607),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7959_ (.CLK(clknet_leaf_20_clk),
    .D(net645),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7960_ (.CLK(clknet_leaf_5_clk),
    .D(net665),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7961_ (.CLK(clknet_leaf_4_clk),
    .D(net669),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7962_ (.CLK(clknet_leaf_46_clk),
    .D(net631),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7963_ (.CLK(clknet_leaf_50_clk),
    .D(net686),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7964_ (.CLK(clknet_leaf_24_clk),
    .D(net759),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7965_ (.CLK(clknet_leaf_53_clk),
    .D(net694),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7966_ (.CLK(clknet_leaf_63_clk),
    .D(net563),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7967_ (.CLK(clknet_leaf_65_clk),
    .D(net633),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7968_ (.CLK(clknet_leaf_69_clk),
    .D(net559),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7969_ (.CLK(clknet_leaf_64_clk),
    .D(net720),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7970_ (.CLK(clknet_leaf_69_clk),
    .D(net641),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7971_ (.CLK(clknet_leaf_66_clk),
    .D(net621),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7972_ (.CLK(clknet_leaf_65_clk),
    .D(net639),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7973_ (.CLK(clknet_leaf_65_clk),
    .D(net579),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7974_ (.CLK(clknet_leaf_72_clk),
    .D(net561),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7975_ (.CLK(clknet_leaf_69_clk),
    .D(net591),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7976_ (.CLK(clknet_leaf_49_clk),
    .D(net643),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7977_ (.CLK(clknet_leaf_68_clk),
    .D(net571),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7978_ (.CLK(clknet_leaf_49_clk),
    .D(_0855_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7979_ (.CLK(clknet_leaf_51_clk),
    .D(_0856_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7980_ (.CLK(clknet_leaf_72_clk),
    .D(_0857_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7981_ (.CLK(clknet_leaf_18_clk),
    .D(_0858_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7982_ (.CLK(clknet_leaf_14_clk),
    .D(_0859_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7983_ (.CLK(clknet_leaf_18_clk),
    .D(_0860_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7984_ (.CLK(clknet_leaf_19_clk),
    .D(_0861_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7985_ (.CLK(clknet_leaf_18_clk),
    .D(_0862_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7986_ (.CLK(clknet_leaf_18_clk),
    .D(_0863_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7987_ (.CLK(clknet_leaf_14_clk),
    .D(_0864_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7988_ (.CLK(clknet_leaf_19_clk),
    .D(_0865_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7989_ (.CLK(clknet_leaf_4_clk),
    .D(_0866_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7990_ (.CLK(clknet_leaf_14_clk),
    .D(_0867_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7991_ (.CLK(clknet_leaf_49_clk),
    .D(_0868_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7992_ (.CLK(clknet_leaf_19_clk),
    .D(_0869_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7993_ (.CLK(clknet_leaf_18_clk),
    .D(_0870_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7994_ (.CLK(clknet_leaf_44_clk),
    .D(_0871_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7995_ (.CLK(clknet_leaf_52_clk),
    .D(_0872_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7996_ (.CLK(clknet_leaf_24_clk),
    .D(_0873_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7997_ (.CLK(clknet_leaf_51_clk),
    .D(_0874_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7998_ (.CLK(clknet_leaf_63_clk),
    .D(_0875_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7999_ (.CLK(clknet_leaf_65_clk),
    .D(_0876_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8000_ (.CLK(clknet_leaf_75_clk),
    .D(_0877_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8001_ (.CLK(clknet_leaf_64_clk),
    .D(_0878_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8002_ (.CLK(clknet_leaf_69_clk),
    .D(_0879_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8003_ (.CLK(clknet_leaf_64_clk),
    .D(_0880_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8004_ (.CLK(clknet_leaf_65_clk),
    .D(_0881_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8005_ (.CLK(clknet_leaf_65_clk),
    .D(_0882_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8006_ (.CLK(clknet_leaf_72_clk),
    .D(_0883_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8007_ (.CLK(clknet_leaf_69_clk),
    .D(_0884_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8008_ (.CLK(clknet_leaf_49_clk),
    .D(_0885_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8009_ (.CLK(clknet_leaf_66_clk),
    .D(_0886_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8010_ (.CLK(clknet_leaf_12_clk),
    .D(_0887_),
    .Q(\U_DATAPATH.U_EX_MEM.i_funct3_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8011_ (.CLK(clknet_leaf_28_clk),
    .D(_0888_),
    .Q(\U_DATAPATH.U_EX_MEM.i_funct3_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8012_ (.CLK(clknet_leaf_79_clk),
    .D(_0889_),
    .Q(\U_DATAPATH.U_EX_MEM.i_funct3_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8013_ (.CLK(net512),
    .D(_0032_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8014_ (.CLK(net513),
    .D(_0043_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8015_ (.CLK(net514),
    .D(_0054_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8016_ (.CLK(net515),
    .D(_0057_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8017_ (.CLK(net516),
    .D(_0058_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8018_ (.CLK(net517),
    .D(_0059_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8019_ (.CLK(net518),
    .D(_0060_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8020_ (.CLK(net519),
    .D(_0061_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8021_ (.CLK(net520),
    .D(_0062_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8022_ (.CLK(net521),
    .D(_0063_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8023_ (.CLK(net522),
    .D(_0033_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8024_ (.CLK(net523),
    .D(_0034_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8025_ (.CLK(net524),
    .D(_0035_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8026_ (.CLK(net525),
    .D(_0036_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8027_ (.CLK(net526),
    .D(_0037_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8028_ (.CLK(net527),
    .D(_0038_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8029_ (.CLK(net528),
    .D(_0039_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8030_ (.CLK(net529),
    .D(_0040_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8031_ (.CLK(net530),
    .D(_0041_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8032_ (.CLK(net531),
    .D(_0042_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8033_ (.CLK(net532),
    .D(_0044_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8034_ (.CLK(net533),
    .D(_0045_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8035_ (.CLK(net534),
    .D(_0046_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8036_ (.CLK(net535),
    .D(_0047_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8037_ (.CLK(net536),
    .D(_0048_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8038_ (.CLK(net537),
    .D(_0049_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8039_ (.CLK(net538),
    .D(_0050_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8040_ (.CLK(net539),
    .D(_0051_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8041_ (.CLK(net540),
    .D(_0052_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8042_ (.CLK(net541),
    .D(_0053_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8043_ (.CLK(net542),
    .D(_0055_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8044_ (.CLK(net543),
    .D(_0056_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8045_ (.CLK(clknet_leaf_36_clk),
    .D(net811),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8046_ (.CLK(clknet_leaf_36_clk),
    .D(net874),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8047_ (.CLK(clknet_leaf_40_clk),
    .D(net978),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8048_ (.CLK(clknet_leaf_34_clk),
    .D(net1148),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8049_ (.CLK(clknet_leaf_12_clk),
    .D(net1276),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8050_ (.CLK(clknet_leaf_26_clk),
    .D(net1557),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8051_ (.CLK(clknet_leaf_40_clk),
    .D(net1198),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8052_ (.CLK(clknet_leaf_48_clk),
    .D(net1723),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8053_ (.CLK(clknet_leaf_14_clk),
    .D(net1140),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8054_ (.CLK(clknet_leaf_34_clk),
    .D(net988),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8055_ (.CLK(clknet_leaf_24_clk),
    .D(net1052),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8056_ (.CLK(clknet_leaf_45_clk),
    .D(net1124),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8057_ (.CLK(clknet_leaf_28_clk),
    .D(net1322),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8058_ (.CLK(clknet_leaf_43_clk),
    .D(net1150),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8059_ (.CLK(clknet_leaf_21_clk),
    .D(net1214),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8060_ (.CLK(clknet_leaf_13_clk),
    .D(net1294),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8061_ (.CLK(clknet_leaf_45_clk),
    .D(net1182),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8062_ (.CLK(clknet_leaf_76_clk),
    .D(net906),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8063_ (.CLK(clknet_leaf_32_clk),
    .D(net1146),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8064_ (.CLK(clknet_leaf_20_clk),
    .D(net1068),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8065_ (.CLK(clknet_leaf_55_clk),
    .D(net1314),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8066_ (.CLK(clknet_leaf_60_clk),
    .D(net1246),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8067_ (.CLK(clknet_leaf_46_clk),
    .D(net1414),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8068_ (.CLK(clknet_leaf_61_clk),
    .D(net1727),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8069_ (.CLK(clknet_leaf_34_clk),
    .D(net1751),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8070_ (.CLK(clknet_leaf_62_clk),
    .D(net1190),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8071_ (.CLK(clknet_leaf_61_clk),
    .D(net1523),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8072_ (.CLK(clknet_leaf_42_clk),
    .D(net900),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8073_ (.CLK(clknet_leaf_54_clk),
    .D(net1184),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8074_ (.CLK(clknet_leaf_75_clk),
    .D(net1252),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8075_ (.CLK(clknet_leaf_30_clk),
    .D(net1340),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8076_ (.CLK(clknet_leaf_59_clk),
    .D(net893),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8077_ (.CLK(clknet_leaf_37_clk),
    .D(net1799),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8078_ (.CLK(clknet_leaf_36_clk),
    .D(net1803),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8079_ (.CLK(clknet_leaf_37_clk),
    .D(net2094),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8080_ (.CLK(clknet_leaf_35_clk),
    .D(net1825),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8081_ (.CLK(clknet_leaf_27_clk),
    .D(net1801),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8082_ (.CLK(clknet_leaf_26_clk),
    .D(net1894),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8083_ (.CLK(clknet_leaf_41_clk),
    .D(net1841),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8084_ (.CLK(clknet_leaf_23_clk),
    .D(net1831),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8085_ (.CLK(clknet_leaf_25_clk),
    .D(net1917),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8086_ (.CLK(clknet_leaf_34_clk),
    .D(net1938),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8087_ (.CLK(clknet_leaf_23_clk),
    .D(net1942),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8088_ (.CLK(clknet_leaf_57_clk),
    .D(net1877),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8089_ (.CLK(clknet_leaf_28_clk),
    .D(net1951),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8090_ (.CLK(clknet_leaf_42_clk),
    .D(net1747),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8091_ (.CLK(clknet_leaf_21_clk),
    .D(net1839),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8092_ (.CLK(clknet_leaf_26_clk),
    .D(net1813),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8093_ (.CLK(clknet_leaf_44_clk),
    .D(net1892),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8094_ (.CLK(clknet_leaf_76_clk),
    .D(net1867),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8095_ (.CLK(clknet_leaf_32_clk),
    .D(net1852),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8096_ (.CLK(clknet_leaf_50_clk),
    .D(net1731),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8097_ (.CLK(clknet_leaf_62_clk),
    .D(net1835),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8098_ (.CLK(clknet_leaf_60_clk),
    .D(net1847),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8099_ (.CLK(clknet_leaf_46_clk),
    .D(net1964),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8100_ (.CLK(clknet_leaf_60_clk),
    .D(net1896),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8101_ (.CLK(clknet_leaf_30_clk),
    .D(net1782),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8102_ (.CLK(clknet_leaf_61_clk),
    .D(net1911),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8103_ (.CLK(clknet_leaf_60_clk),
    .D(net1930),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8104_ (.CLK(clknet_leaf_41_clk),
    .D(net1909),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8105_ (.CLK(clknet_leaf_53_clk),
    .D(net1898),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8106_ (.CLK(clknet_leaf_55_clk),
    .D(net1786),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8107_ (.CLK(clknet_leaf_29_clk),
    .D(net1907),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8108_ (.CLK(clknet_leaf_43_clk),
    .D(net1769),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8109_ (.CLK(clknet_leaf_37_clk),
    .D(net806),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8110_ (.CLK(clknet_leaf_36_clk),
    .D(net1457),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8111_ (.CLK(clknet_leaf_37_clk),
    .D(net795),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8112_ (.CLK(clknet_leaf_35_clk),
    .D(net1072),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8113_ (.CLK(clknet_leaf_27_clk),
    .D(net1505),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8114_ (.CLK(clknet_leaf_26_clk),
    .D(net1076),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8115_ (.CLK(clknet_leaf_41_clk),
    .D(net1204),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8116_ (.CLK(clknet_leaf_23_clk),
    .D(net1445),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8117_ (.CLK(clknet_leaf_26_clk),
    .D(net1188),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8118_ (.CLK(clknet_leaf_34_clk),
    .D(net1174),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8119_ (.CLK(clknet_leaf_24_clk),
    .D(net1679),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8120_ (.CLK(clknet_leaf_57_clk),
    .D(net1020),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8121_ (.CLK(clknet_leaf_28_clk),
    .D(net1587),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8122_ (.CLK(clknet_leaf_42_clk),
    .D(net1128),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8123_ (.CLK(clknet_leaf_21_clk),
    .D(net1372),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8124_ (.CLK(clknet_leaf_27_clk),
    .D(net1036),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8125_ (.CLK(clknet_leaf_46_clk),
    .D(net1499),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8126_ (.CLK(clknet_leaf_54_clk),
    .D(net1222),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8127_ (.CLK(clknet_leaf_33_clk),
    .D(net1485),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8128_ (.CLK(clknet_leaf_51_clk),
    .D(net1008),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8129_ (.CLK(clknet_leaf_55_clk),
    .D(net1208),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8130_ (.CLK(clknet_leaf_60_clk),
    .D(net1567),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8131_ (.CLK(clknet_leaf_46_clk),
    .D(net1589),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8132_ (.CLK(clknet_leaf_61_clk),
    .D(net1310),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8133_ (.CLK(clknet_leaf_30_clk),
    .D(net980),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8134_ (.CLK(clknet_leaf_62_clk),
    .D(net1569),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8135_ (.CLK(clknet_leaf_60_clk),
    .D(net1753),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8136_ (.CLK(clknet_leaf_41_clk),
    .D(net1455),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8137_ (.CLK(clknet_leaf_53_clk),
    .D(net982),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8138_ (.CLK(clknet_leaf_55_clk),
    .D(net1491),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8139_ (.CLK(clknet_leaf_29_clk),
    .D(net1122),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8140_ (.CLK(clknet_leaf_43_clk),
    .D(net1702),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8141_ (.CLK(clknet_leaf_38_clk),
    .D(net912),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8142_ (.CLK(clknet_leaf_38_clk),
    .D(net1296),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8143_ (.CLK(clknet_leaf_39_clk),
    .D(net1200),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8144_ (.CLK(clknet_leaf_38_clk),
    .D(net868),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8145_ (.CLK(clknet_leaf_28_clk),
    .D(net1437),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8146_ (.CLK(clknet_leaf_25_clk),
    .D(net1336),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8147_ (.CLK(clknet_leaf_39_clk),
    .D(net1010),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8148_ (.CLK(clknet_leaf_23_clk),
    .D(net1406),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8149_ (.CLK(clknet_leaf_23_clk),
    .D(net1206),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8150_ (.CLK(clknet_leaf_33_clk),
    .D(net1238),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8151_ (.CLK(clknet_leaf_25_clk),
    .D(net1384),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8152_ (.CLK(clknet_leaf_56_clk),
    .D(net1186),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8153_ (.CLK(clknet_leaf_29_clk),
    .D(net1394),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8154_ (.CLK(clknet_leaf_44_clk),
    .D(net1593),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8155_ (.CLK(clknet_leaf_48_clk),
    .D(net1577),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8156_ (.CLK(clknet_leaf_25_clk),
    .D(net1386),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8157_ (.CLK(clknet_leaf_49_clk),
    .D(net1439),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8158_ (.CLK(clknet_leaf_52_clk),
    .D(net1416),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8159_ (.CLK(clknet_leaf_24_clk),
    .D(net1278),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8160_ (.CLK(clknet_leaf_50_clk),
    .D(net928),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8161_ (.CLK(clknet_leaf_54_clk),
    .D(net1541),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8162_ (.CLK(clknet_leaf_58_clk),
    .D(net1757),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8163_ (.CLK(clknet_leaf_47_clk),
    .D(net1274),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8164_ (.CLK(clknet_leaf_62_clk),
    .D(net1461),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8165_ (.CLK(clknet_leaf_30_clk),
    .D(net1344),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8166_ (.CLK(clknet_leaf_56_clk),
    .D(net1398),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8167_ (.CLK(clknet_leaf_60_clk),
    .D(net1561),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8168_ (.CLK(clknet_leaf_40_clk),
    .D(net1046),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8169_ (.CLK(clknet_leaf_53_clk),
    .D(net1162),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8170_ (.CLK(clknet_leaf_54_clk),
    .D(net1212),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8171_ (.CLK(clknet_leaf_29_clk),
    .D(net1006),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8172_ (.CLK(clknet_leaf_44_clk),
    .D(net1192),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8173_ (.CLK(clknet_leaf_38_clk),
    .D(net1932),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8174_ (.CLK(clknet_leaf_36_clk),
    .D(net1819),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8175_ (.CLK(clknet_leaf_40_clk),
    .D(net1685),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8176_ (.CLK(clknet_leaf_33_clk),
    .D(net2103),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8177_ (.CLK(clknet_leaf_28_clk),
    .D(net1981),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8178_ (.CLK(clknet_leaf_24_clk),
    .D(net1763),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8179_ (.CLK(clknet_leaf_40_clk),
    .D(net1871),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8180_ (.CLK(clknet_leaf_48_clk),
    .D(net1900),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8181_ (.CLK(clknet_leaf_23_clk),
    .D(net1949),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8182_ (.CLK(clknet_leaf_35_clk),
    .D(net1710),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8183_ (.CLK(clknet_leaf_25_clk),
    .D(net1773),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8184_ (.CLK(clknet_leaf_57_clk),
    .D(net1859),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8185_ (.CLK(clknet_leaf_29_clk),
    .D(net1927),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8186_ (.CLK(clknet_leaf_44_clk),
    .D(net1861),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8187_ (.CLK(clknet_leaf_23_clk),
    .D(net1957),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8188_ (.CLK(clknet_leaf_25_clk),
    .D(net1623),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8189_ (.CLK(clknet_leaf_45_clk),
    .D(net1663),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8190_ (.CLK(clknet_leaf_54_clk),
    .D(net1903),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8191_ (.CLK(clknet_leaf_32_clk),
    .D(net1821),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8192_ (.CLK(clknet_leaf_49_clk),
    .D(net1735),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8193_ (.CLK(clknet_leaf_56_clk),
    .D(net1884),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8194_ (.CLK(clknet_leaf_59_clk),
    .D(net1777),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8195_ (.CLK(clknet_leaf_46_clk),
    .D(net1966),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8196_ (.CLK(clknet_leaf_60_clk),
    .D(net1923),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8197_ (.CLK(clknet_leaf_33_clk),
    .D(net1925),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8198_ (.CLK(clknet_leaf_62_clk),
    .D(net1915),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8199_ (.CLK(clknet_leaf_60_clk),
    .D(net1913),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8200_ (.CLK(clknet_leaf_42_clk),
    .D(net1765),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8201_ (.CLK(clknet_leaf_56_clk),
    .D(net1890),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8202_ (.CLK(clknet_leaf_54_clk),
    .D(net1979),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8203_ (.CLK(clknet_leaf_30_clk),
    .D(net1796),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8204_ (.CLK(clknet_leaf_43_clk),
    .D(net1706),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8205_ (.CLK(clknet_leaf_37_clk),
    .D(net785),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8206_ (.CLK(clknet_leaf_38_clk),
    .D(net1809),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8207_ (.CLK(clknet_leaf_37_clk),
    .D(net798),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8208_ (.CLK(clknet_leaf_33_clk),
    .D(net1471),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8209_ (.CLK(clknet_leaf_28_clk),
    .D(net1388),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8210_ (.CLK(clknet_leaf_26_clk),
    .D(net1090),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8211_ (.CLK(clknet_leaf_41_clk),
    .D(net1260),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8212_ (.CLK(clknet_leaf_23_clk),
    .D(net1533),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8213_ (.CLK(clknet_leaf_26_clk),
    .D(net1429),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8214_ (.CLK(clknet_leaf_34_clk),
    .D(net1158),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8215_ (.CLK(clknet_leaf_23_clk),
    .D(net1453),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8216_ (.CLK(clknet_leaf_57_clk),
    .D(net1509),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8217_ (.CLK(clknet_leaf_28_clk),
    .D(net1549),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8218_ (.CLK(clknet_leaf_43_clk),
    .D(net1376),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8219_ (.CLK(clknet_leaf_21_clk),
    .D(net1080),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8220_ (.CLK(clknet_leaf_27_clk),
    .D(net1242),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8221_ (.CLK(clknet_leaf_45_clk),
    .D(net964),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8222_ (.CLK(clknet_leaf_76_clk),
    .D(net908),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8223_ (.CLK(clknet_leaf_31_clk),
    .D(net1493),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8224_ (.CLK(clknet_leaf_20_clk),
    .D(net994),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8225_ (.CLK(clknet_leaf_55_clk),
    .D(net1423),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8226_ (.CLK(clknet_leaf_60_clk),
    .D(net1334),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8227_ (.CLK(clknet_leaf_46_clk),
    .D(net1627),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8228_ (.CLK(clknet_leaf_61_clk),
    .D(net1575),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8229_ (.CLK(clknet_leaf_30_clk),
    .D(net974),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8230_ (.CLK(clknet_leaf_56_clk),
    .D(net1689),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8231_ (.CLK(clknet_leaf_60_clk),
    .D(net1537),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8232_ (.CLK(clknet_leaf_41_clk),
    .D(net1435),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8233_ (.CLK(clknet_leaf_52_clk),
    .D(net943),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8234_ (.CLK(clknet_leaf_75_clk),
    .D(net1270),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8235_ (.CLK(clknet_leaf_28_clk),
    .D(net1515),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8236_ (.CLK(clknet_leaf_43_clk),
    .D(net986),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8237_ (.CLK(clknet_leaf_37_clk),
    .D(net941),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8238_ (.CLK(clknet_leaf_38_clk),
    .D(net1968),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8239_ (.CLK(clknet_leaf_37_clk),
    .D(net787),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8240_ (.CLK(clknet_leaf_33_clk),
    .D(net1316),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8241_ (.CLK(clknet_leaf_27_clk),
    .D(net1306),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8242_ (.CLK(clknet_leaf_13_clk),
    .D(net1390),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8243_ (.CLK(clknet_leaf_41_clk),
    .D(net1364),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8244_ (.CLK(clknet_leaf_23_clk),
    .D(net1244),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8245_ (.CLK(clknet_leaf_26_clk),
    .D(net1360),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8246_ (.CLK(clknet_leaf_34_clk),
    .D(net1487),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8247_ (.CLK(clknet_leaf_23_clk),
    .D(net1525),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8248_ (.CLK(clknet_leaf_57_clk),
    .D(net1298),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8249_ (.CLK(clknet_leaf_28_clk),
    .D(net1142),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8250_ (.CLK(clknet_leaf_43_clk),
    .D(net1110),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8251_ (.CLK(clknet_leaf_21_clk),
    .D(net1312),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8252_ (.CLK(clknet_leaf_27_clk),
    .D(net1302),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8253_ (.CLK(clknet_leaf_45_clk),
    .D(net1144),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8254_ (.CLK(clknet_leaf_76_clk),
    .D(net1226),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8255_ (.CLK(clknet_leaf_31_clk),
    .D(net1531),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8256_ (.CLK(clknet_leaf_20_clk),
    .D(net1028),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8257_ (.CLK(clknet_leaf_55_clk),
    .D(net1082),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8258_ (.CLK(clknet_leaf_60_clk),
    .D(net1138),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8259_ (.CLK(clknet_leaf_46_clk),
    .D(net1649),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8260_ (.CLK(clknet_leaf_61_clk),
    .D(net1164),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8261_ (.CLK(clknet_leaf_29_clk),
    .D(net918),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8262_ (.CLK(clknet_leaf_62_clk),
    .D(net1272),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8263_ (.CLK(clknet_leaf_60_clk),
    .D(net1092),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8264_ (.CLK(clknet_leaf_42_clk),
    .D(net945),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8265_ (.CLK(clknet_leaf_53_clk),
    .D(net992),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8266_ (.CLK(clknet_leaf_75_clk),
    .D(net1402),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8267_ (.CLK(clknet_leaf_29_clk),
    .D(net1332),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8268_ (.CLK(clknet_leaf_59_clk),
    .D(net933),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ));
 sky130_fd_sc_hd__dfstp_1 _8269_ (.CLK(clknet_leaf_73_clk),
    .D(_1114_),
    .SET_B(_0163_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8270_ (.CLK(clknet_leaf_17_clk),
    .D(_1115_),
    .RESET_B(_0164_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8271_ (.CLK(clknet_leaf_16_clk),
    .D(_1116_),
    .RESET_B(_0165_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8272_ (.CLK(clknet_leaf_7_clk),
    .D(net1994),
    .RESET_B(_0166_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8273_ (.CLK(clknet_leaf_16_clk),
    .D(_1118_),
    .RESET_B(_0167_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8274_ (.CLK(clknet_leaf_16_clk),
    .D(_1119_),
    .RESET_B(_0168_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8275_ (.CLK(clknet_leaf_16_clk),
    .D(_1120_),
    .RESET_B(_0169_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8276_ (.CLK(clknet_leaf_15_clk),
    .D(net2014),
    .RESET_B(_0170_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8277_ (.CLK(clknet_leaf_6_clk),
    .D(net2045),
    .RESET_B(_0171_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8278_ (.CLK(clknet_leaf_6_clk),
    .D(_1123_),
    .RESET_B(_0172_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8279_ (.CLK(clknet_leaf_7_clk),
    .D(_1124_),
    .RESET_B(_0173_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8280_ (.CLK(clknet_leaf_5_clk),
    .D(_1125_),
    .RESET_B(_0174_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8281_ (.CLK(clknet_leaf_5_clk),
    .D(_1126_),
    .RESET_B(_0175_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8282_ (.CLK(clknet_leaf_5_clk),
    .D(_1127_),
    .RESET_B(_0176_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8283_ (.CLK(clknet_leaf_48_clk),
    .D(_1128_),
    .RESET_B(_0177_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8284_ (.CLK(clknet_leaf_48_clk),
    .D(_1129_),
    .RESET_B(_0178_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8285_ (.CLK(clknet_leaf_49_clk),
    .D(_1130_),
    .RESET_B(_0179_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8286_ (.CLK(clknet_leaf_53_clk),
    .D(_1131_),
    .RESET_B(_0180_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[19] ));
 sky130_fd_sc_hd__dfrtp_1 _8287_ (.CLK(clknet_leaf_75_clk),
    .D(net2065),
    .RESET_B(_0181_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[20] ));
 sky130_fd_sc_hd__dfrtp_1 _8288_ (.CLK(clknet_leaf_63_clk),
    .D(_1133_),
    .RESET_B(_0182_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8289_ (.CLK(clknet_leaf_63_clk),
    .D(_1134_),
    .RESET_B(_0183_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8290_ (.CLK(clknet_leaf_64_clk),
    .D(net2022),
    .RESET_B(_0184_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8291_ (.CLK(clknet_leaf_68_clk),
    .D(_1136_),
    .RESET_B(_0185_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8292_ (.CLK(clknet_leaf_67_clk),
    .D(_1137_),
    .RESET_B(_0186_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[25] ));
 sky130_fd_sc_hd__dfrtp_1 _8293_ (.CLK(clknet_leaf_68_clk),
    .D(_1138_),
    .RESET_B(_0187_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8294_ (.CLK(clknet_leaf_68_clk),
    .D(_1139_),
    .RESET_B(_0188_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[27] ));
 sky130_fd_sc_hd__dfrtp_1 _8295_ (.CLK(clknet_leaf_71_clk),
    .D(_1140_),
    .RESET_B(_0189_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[28] ));
 sky130_fd_sc_hd__dfrtp_1 _8296_ (.CLK(clknet_leaf_71_clk),
    .D(_1141_),
    .RESET_B(_0190_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[29] ));
 sky130_fd_sc_hd__dfrtp_1 _8297_ (.CLK(clknet_leaf_71_clk),
    .D(_1142_),
    .RESET_B(_0191_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[30] ));
 sky130_fd_sc_hd__dfrtp_1 _8298_ (.CLK(clknet_leaf_71_clk),
    .D(_1143_),
    .RESET_B(_0192_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8299_ (.CLK(clknet_leaf_38_clk),
    .D(net1953),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8300_ (.CLK(clknet_leaf_35_clk),
    .D(net2087),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8301_ (.CLK(clknet_leaf_40_clk),
    .D(net1741),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8302_ (.CLK(clknet_leaf_34_clk),
    .D(net1629),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8303_ (.CLK(clknet_leaf_12_clk),
    .D(net1637),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8304_ (.CLK(clknet_leaf_13_clk),
    .D(net2128),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8305_ (.CLK(clknet_leaf_40_clk),
    .D(net1745),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8306_ (.CLK(clknet_leaf_23_clk),
    .D(net1771),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8307_ (.CLK(clknet_leaf_14_clk),
    .D(net1886),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8308_ (.CLK(clknet_leaf_34_clk),
    .D(net1667),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8309_ (.CLK(clknet_leaf_25_clk),
    .D(net1759),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8310_ (.CLK(clknet_leaf_45_clk),
    .D(net1704),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8311_ (.CLK(clknet_leaf_28_clk),
    .D(net1921),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8312_ (.CLK(clknet_leaf_43_clk),
    .D(net1761),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8313_ (.CLK(clknet_leaf_21_clk),
    .D(net1837),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8314_ (.CLK(clknet_leaf_13_clk),
    .D(net1849),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8315_ (.CLK(clknet_leaf_45_clk),
    .D(net1697),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8316_ (.CLK(clknet_leaf_76_clk),
    .D(net1545),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8317_ (.CLK(clknet_leaf_32_clk),
    .D(net1829),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8318_ (.CLK(clknet_leaf_20_clk),
    .D(net1659),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8319_ (.CLK(clknet_leaf_55_clk),
    .D(net1779),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8320_ (.CLK(clknet_leaf_58_clk),
    .D(net1749),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8321_ (.CLK(clknet_leaf_46_clk),
    .D(net1940),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8322_ (.CLK(clknet_leaf_61_clk),
    .D(net1784),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8323_ (.CLK(clknet_leaf_30_clk),
    .D(net1811),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8324_ (.CLK(clknet_leaf_62_clk),
    .D(net1794),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8325_ (.CLK(clknet_leaf_61_clk),
    .D(net1712),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8326_ (.CLK(clknet_leaf_42_clk),
    .D(net1603),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8327_ (.CLK(clknet_leaf_54_clk),
    .D(net1792),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8328_ (.CLK(clknet_leaf_75_clk),
    .D(net1823),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8329_ (.CLK(clknet_leaf_29_clk),
    .D(net1857),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8330_ (.CLK(clknet_leaf_59_clk),
    .D(net1529),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8331_ (.CLK(clknet_leaf_36_clk),
    .D(net2082),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8332_ (.CLK(clknet_leaf_36_clk),
    .D(net1565),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8333_ (.CLK(clknet_leaf_41_clk),
    .D(net1657),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8334_ (.CLK(clknet_leaf_35_clk),
    .D(net1755),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8335_ (.CLK(clknet_leaf_28_clk),
    .D(net1976),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8336_ (.CLK(clknet_leaf_14_clk),
    .D(net2115),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8337_ (.CLK(clknet_leaf_41_clk),
    .D(net1665),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8338_ (.CLK(clknet_leaf_48_clk),
    .D(net1739),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8339_ (.CLK(clknet_leaf_22_clk),
    .D(net1717),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8340_ (.CLK(clknet_leaf_34_clk),
    .D(net1790),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8341_ (.CLK(clknet_leaf_24_clk),
    .D(net1843),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8342_ (.CLK(clknet_leaf_44_clk),
    .D(net1959),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8343_ (.CLK(clknet_leaf_28_clk),
    .D(net1970),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8344_ (.CLK(clknet_leaf_43_clk),
    .D(net1833),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8345_ (.CLK(clknet_leaf_21_clk),
    .D(net1873),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8346_ (.CLK(clknet_leaf_26_clk),
    .D(net1845),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8347_ (.CLK(clknet_leaf_44_clk),
    .D(net1882),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8348_ (.CLK(clknet_leaf_75_clk),
    .D(net1919),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8349_ (.CLK(clknet_leaf_32_clk),
    .D(net1647),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8350_ (.CLK(clknet_leaf_20_clk),
    .D(net1767),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8351_ (.CLK(clknet_leaf_62_clk),
    .D(net1807),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8352_ (.CLK(clknet_leaf_59_clk),
    .D(net1617),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8353_ (.CLK(clknet_leaf_46_clk),
    .D(net1936),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8354_ (.CLK(clknet_leaf_61_clk),
    .D(net1863),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8355_ (.CLK(clknet_leaf_30_clk),
    .D(net1817),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8356_ (.CLK(clknet_leaf_62_clk),
    .D(net1788),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8357_ (.CLK(clknet_leaf_61_clk),
    .D(net1962),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8358_ (.CLK(clknet_leaf_42_clk),
    .D(net1443),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8359_ (.CLK(clknet_leaf_54_clk),
    .D(net1854),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8360_ (.CLK(clknet_leaf_75_clk),
    .D(net1905),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8361_ (.CLK(clknet_leaf_29_clk),
    .D(net1865),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8362_ (.CLK(clknet_leaf_59_clk),
    .D(net1563),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8363_ (.CLK(clknet_leaf_2_clk),
    .D(_1208_),
    .Q(\U_DATAPATH.U_EX_MEM.i_result_src_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8364_ (.CLK(clknet_leaf_78_clk),
    .D(net2207),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8365_ (.CLK(clknet_leaf_78_clk),
    .D(_1210_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8366_ (.CLK(clknet_leaf_78_clk),
    .D(_1211_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8367_ (.CLK(clknet_leaf_78_clk),
    .D(_1212_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8368_ (.CLK(clknet_leaf_37_clk),
    .D(net1591),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8369_ (.CLK(clknet_leaf_36_clk),
    .D(net1553),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8370_ (.CLK(clknet_leaf_41_clk),
    .D(net1154),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8371_ (.CLK(clknet_leaf_35_clk),
    .D(net1290),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8372_ (.CLK(clknet_leaf_12_clk),
    .D(net1104),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8373_ (.CLK(clknet_leaf_26_clk),
    .D(net1404),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8374_ (.CLK(clknet_leaf_41_clk),
    .D(net1677),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8375_ (.CLK(clknet_leaf_47_clk),
    .D(net1210),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8376_ (.CLK(clknet_leaf_26_clk),
    .D(net1599),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8377_ (.CLK(clknet_leaf_34_clk),
    .D(net1427),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8378_ (.CLK(clknet_leaf_24_clk),
    .D(net1609),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8379_ (.CLK(clknet_leaf_44_clk),
    .D(net1708),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8380_ (.CLK(clknet_leaf_28_clk),
    .D(net1643),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8381_ (.CLK(clknet_leaf_43_clk),
    .D(net1378),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8382_ (.CLK(clknet_leaf_22_clk),
    .D(net1266),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8383_ (.CLK(clknet_leaf_27_clk),
    .D(net1683),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8384_ (.CLK(clknet_leaf_44_clk),
    .D(net1483),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8385_ (.CLK(clknet_leaf_75_clk),
    .D(net1631),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8386_ (.CLK(clknet_leaf_32_clk),
    .D(net1721),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8387_ (.CLK(clknet_leaf_20_clk),
    .D(net1342),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8388_ (.CLK(clknet_leaf_62_clk),
    .D(net1473),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8389_ (.CLK(clknet_leaf_59_clk),
    .D(net1088),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8390_ (.CLK(clknet_leaf_39_clk),
    .D(net1451),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8391_ (.CLK(clknet_leaf_61_clk),
    .D(net1595),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8392_ (.CLK(clknet_leaf_30_clk),
    .D(net1380),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8393_ (.CLK(clknet_leaf_62_clk),
    .D(net1601),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8394_ (.CLK(clknet_leaf_61_clk),
    .D(net1607),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8395_ (.CLK(clknet_leaf_42_clk),
    .D(net1054),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8396_ (.CLK(clknet_leaf_53_clk),
    .D(net1421),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8397_ (.CLK(clknet_leaf_75_clk),
    .D(net1539),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8398_ (.CLK(clknet_leaf_30_clk),
    .D(net1733),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8399_ (.CLK(clknet_leaf_59_clk),
    .D(net1513),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8400_ (.CLK(clknet_leaf_80_clk),
    .D(_1245_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8401_ (.CLK(clknet_leaf_70_clk),
    .D(_1246_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8402_ (.CLK(clknet_leaf_73_clk),
    .D(_1247_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8403_ (.CLK(clknet_leaf_80_clk),
    .D(net2003),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8404_ (.CLK(clknet_leaf_74_clk),
    .D(_1249_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8405_ (.CLK(clknet_leaf_74_clk),
    .D(net1974),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8406_ (.CLK(clknet_leaf_74_clk),
    .D(net2020),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8407_ (.CLK(clknet_leaf_74_clk),
    .D(_1252_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8408_ (.CLK(clknet_leaf_74_clk),
    .D(_1253_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8409_ (.CLK(clknet_leaf_75_clk),
    .D(_1254_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8410_ (.CLK(clknet_leaf_75_clk),
    .D(_1255_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8411_ (.CLK(clknet_leaf_75_clk),
    .D(_1256_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8412_ (.CLK(clknet_leaf_51_clk),
    .D(_1257_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8413_ (.CLK(clknet_leaf_50_clk),
    .D(net1947),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8414_ (.CLK(clknet_leaf_51_clk),
    .D(_1259_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8415_ (.CLK(clknet_leaf_51_clk),
    .D(_1260_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8416_ (.CLK(clknet_leaf_20_clk),
    .D(_1261_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8417_ (.CLK(clknet_leaf_4_clk),
    .D(_1262_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8418_ (.CLK(clknet_leaf_4_clk),
    .D(_1263_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8419_ (.CLK(clknet_leaf_4_clk),
    .D(net1700),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8420_ (.CLK(clknet_leaf_2_clk),
    .D(_1265_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8421_ (.CLK(clknet_leaf_5_clk),
    .D(_1266_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8422_ (.CLK(clknet_leaf_5_clk),
    .D(_1267_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ));
 sky130_fd_sc_hd__dfxtp_2 _8423_ (.CLK(clknet_leaf_78_clk),
    .D(net1743),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8424_ (.CLK(clknet_leaf_3_clk),
    .D(_1269_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8425_ (.CLK(clknet_leaf_5_clk),
    .D(_1270_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8426_ (.CLK(clknet_leaf_3_clk),
    .D(_1271_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8427_ (.CLK(clknet_leaf_3_clk),
    .D(_1272_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8428_ (.CLK(clknet_leaf_51_clk),
    .D(_1273_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8429_ (.CLK(clknet_leaf_77_clk),
    .D(_1274_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8430_ (.CLK(clknet_leaf_77_clk),
    .D(_1275_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8431_ (.CLK(clknet_leaf_3_clk),
    .D(_1276_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[0] ));
 sky130_fd_sc_hd__ebufn_1 _8439_ (.A(net478),
    .TE_B(_3622_),
    .Z(_0064_));
 sky130_fd_sc_hd__conb_1 _8439__478 (.HI(net478));
 sky130_fd_sc_hd__ebufn_1 _8440_ (.A(net479),
    .TE_B(_3623_),
    .Z(_0065_));
 sky130_fd_sc_hd__conb_1 _8440__479 (.HI(net479));
 sky130_fd_sc_hd__ebufn_1 _8441_ (.A(net473),
    .TE_B(_3624_),
    .Z(_0066_));
 sky130_fd_sc_hd__conb_1 _8441__473 (.LO(net473));
 sky130_fd_sc_hd__ebufn_1 _8442_ (.A(net474),
    .TE_B(_3625_),
    .Z(_0067_));
 sky130_fd_sc_hd__conb_1 _8442__474 (.LO(net474));
 sky130_fd_sc_hd__ebufn_1 _8443_ (.A(net475),
    .TE_B(_3626_),
    .Z(_0068_));
 sky130_fd_sc_hd__conb_1 _8443__475 (.LO(net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__conb_1 core_476 (.LO(net476));
 sky130_fd_sc_hd__conb_1 core_477 (.LO(net477));
 sky130_fd_sc_hd__buf_8 fanout162 (.A(_2647_),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 fanout163 (.A(_2647_),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_8 fanout164 (.A(net166),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_4 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_8 fanout167 (.A(_2522_),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_8 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__buf_6 fanout169 (.A(_2522_),
    .X(net169));
 sky130_fd_sc_hd__buf_6 fanout170 (.A(_2522_),
    .X(net170));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(net173),
    .X(net171));
 sky130_fd_sc_hd__buf_4 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(net2085),
    .X(net173));
 sky130_fd_sc_hd__buf_6 fanout174 (.A(net183),
    .X(net174));
 sky130_fd_sc_hd__buf_4 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__buf_4 fanout176 (.A(net178),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_8 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_8 fanout178 (.A(net183),
    .X(net178));
 sky130_fd_sc_hd__buf_6 fanout179 (.A(net182),
    .X(net179));
 sky130_fd_sc_hd__buf_4 fanout180 (.A(net182),
    .X(net180));
 sky130_fd_sc_hd__buf_4 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__buf_6 fanout182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_8 fanout183 (.A(_1780_),
    .X(net183));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(_1589_),
    .X(net185));
 sky130_fd_sc_hd__buf_4 fanout186 (.A(_1589_),
    .X(net186));
 sky130_fd_sc_hd__buf_2 fanout187 (.A(_1589_),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_8 fanout188 (.A(net190),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_8 fanout190 (.A(_1588_),
    .X(net190));
 sky130_fd_sc_hd__buf_4 fanout191 (.A(net195),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_8 fanout192 (.A(net195),
    .X(net192));
 sky130_fd_sc_hd__buf_4 fanout193 (.A(net195),
    .X(net193));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__buf_4 fanout195 (.A(_1567_),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_8 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_8 fanout197 (.A(net198),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_8 fanout198 (.A(_1556_),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_8 fanout199 (.A(_1555_),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_8 fanout200 (.A(_1555_),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_8 fanout201 (.A(net203),
    .X(net201));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_8 fanout203 (.A(_1540_),
    .X(net203));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(_1539_),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_4 fanout205 (.A(_1539_),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_8 fanout206 (.A(_1539_),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_8 fanout207 (.A(net210),
    .X(net207));
 sky130_fd_sc_hd__buf_2 fanout208 (.A(net210),
    .X(net208));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__buf_2 fanout210 (.A(_1528_),
    .X(net210));
 sky130_fd_sc_hd__buf_4 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__buf_4 fanout212 (.A(net214),
    .X(net212));
 sky130_fd_sc_hd__buf_4 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(_1527_),
    .X(net214));
 sky130_fd_sc_hd__buf_8 fanout215 (.A(_3500_),
    .X(net215));
 sky130_fd_sc_hd__buf_8 fanout216 (.A(_3500_),
    .X(net216));
 sky130_fd_sc_hd__buf_8 fanout217 (.A(_3458_),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_8 fanout218 (.A(_3458_),
    .X(net218));
 sky130_fd_sc_hd__buf_8 fanout219 (.A(_3453_),
    .X(net219));
 sky130_fd_sc_hd__buf_6 fanout220 (.A(_3453_),
    .X(net220));
 sky130_fd_sc_hd__buf_6 fanout221 (.A(_2737_),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_8 fanout222 (.A(net224),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_8 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__buf_6 fanout224 (.A(_2736_),
    .X(net224));
 sky130_fd_sc_hd__buf_6 fanout225 (.A(_2644_),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_8 fanout226 (.A(_2644_),
    .X(net226));
 sky130_fd_sc_hd__buf_6 fanout227 (.A(_2640_),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_8 fanout228 (.A(_2640_),
    .X(net228));
 sky130_fd_sc_hd__buf_6 fanout229 (.A(_2635_),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_8 fanout230 (.A(_2635_),
    .X(net230));
 sky130_fd_sc_hd__buf_8 fanout231 (.A(_2631_),
    .X(net231));
 sky130_fd_sc_hd__buf_6 fanout232 (.A(_2631_),
    .X(net232));
 sky130_fd_sc_hd__buf_8 fanout233 (.A(_2626_),
    .X(net233));
 sky130_fd_sc_hd__buf_6 fanout234 (.A(_2626_),
    .X(net234));
 sky130_fd_sc_hd__buf_6 fanout235 (.A(_2620_),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_8 fanout236 (.A(_2620_),
    .X(net236));
 sky130_fd_sc_hd__buf_8 fanout237 (.A(net238),
    .X(net237));
 sky130_fd_sc_hd__buf_8 fanout238 (.A(_3537_),
    .X(net238));
 sky130_fd_sc_hd__buf_6 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__buf_8 fanout240 (.A(_3536_),
    .X(net240));
 sky130_fd_sc_hd__buf_8 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__buf_8 fanout242 (.A(_3503_),
    .X(net242));
 sky130_fd_sc_hd__buf_6 fanout243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__buf_8 fanout244 (.A(_3502_),
    .X(net244));
 sky130_fd_sc_hd__buf_8 fanout245 (.A(_3498_),
    .X(net245));
 sky130_fd_sc_hd__buf_8 fanout246 (.A(_3498_),
    .X(net246));
 sky130_fd_sc_hd__buf_8 fanout247 (.A(_3496_),
    .X(net247));
 sky130_fd_sc_hd__buf_6 fanout248 (.A(_3496_),
    .X(net248));
 sky130_fd_sc_hd__buf_8 fanout249 (.A(_3461_),
    .X(net249));
 sky130_fd_sc_hd__buf_6 fanout250 (.A(_3461_),
    .X(net250));
 sky130_fd_sc_hd__buf_6 fanout251 (.A(_3460_),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_8 fanout252 (.A(_3460_),
    .X(net252));
 sky130_fd_sc_hd__buf_8 fanout253 (.A(_3456_),
    .X(net253));
 sky130_fd_sc_hd__buf_6 fanout254 (.A(_3456_),
    .X(net254));
 sky130_fd_sc_hd__buf_8 fanout255 (.A(_3451_),
    .X(net255));
 sky130_fd_sc_hd__buf_8 fanout256 (.A(_3451_),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_16 fanout257 (.A(_3414_),
    .X(net257));
 sky130_fd_sc_hd__buf_6 fanout258 (.A(_3414_),
    .X(net258));
 sky130_fd_sc_hd__buf_6 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__buf_8 fanout260 (.A(_2642_),
    .X(net260));
 sky130_fd_sc_hd__buf_6 fanout261 (.A(_2638_),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_8 fanout262 (.A(_2638_),
    .X(net262));
 sky130_fd_sc_hd__buf_6 fanout263 (.A(_2633_),
    .X(net263));
 sky130_fd_sc_hd__buf_6 fanout264 (.A(_2633_),
    .X(net264));
 sky130_fd_sc_hd__buf_8 fanout265 (.A(_2629_),
    .X(net265));
 sky130_fd_sc_hd__buf_8 fanout266 (.A(_2629_),
    .X(net266));
 sky130_fd_sc_hd__buf_8 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__buf_8 fanout268 (.A(_2624_),
    .X(net268));
 sky130_fd_sc_hd__buf_6 fanout269 (.A(_2618_),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_8 fanout270 (.A(_2618_),
    .X(net270));
 sky130_fd_sc_hd__buf_4 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__buf_4 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__buf_2 fanout273 (.A(net291),
    .X(net273));
 sky130_fd_sc_hd__buf_4 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__buf_4 fanout275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_8 fanout276 (.A(net291),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_8 fanout277 (.A(net291),
    .X(net277));
 sky130_fd_sc_hd__buf_2 fanout278 (.A(net291),
    .X(net278));
 sky130_fd_sc_hd__buf_4 fanout279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__buf_4 fanout280 (.A(net283),
    .X(net280));
 sky130_fd_sc_hd__buf_4 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_4 fanout282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 fanout283 (.A(net291),
    .X(net283));
 sky130_fd_sc_hd__buf_4 fanout284 (.A(net286),
    .X(net284));
 sky130_fd_sc_hd__buf_4 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__buf_4 fanout286 (.A(net291),
    .X(net286));
 sky130_fd_sc_hd__buf_4 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 fanout288 (.A(net289),
    .X(net288));
 sky130_fd_sc_hd__buf_4 fanout289 (.A(net291),
    .X(net289));
 sky130_fd_sc_hd__buf_4 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__buf_8 fanout291 (.A(_2076_),
    .X(net291));
 sky130_fd_sc_hd__buf_4 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__buf_4 fanout293 (.A(net295),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_8 fanout294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_8 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__buf_6 fanout296 (.A(_2075_),
    .X(net296));
 sky130_fd_sc_hd__buf_4 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_8 fanout298 (.A(net299),
    .X(net298));
 sky130_fd_sc_hd__buf_6 fanout299 (.A(_2075_),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_8 fanout300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__buf_8 fanout302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_16 fanout303 (.A(_1336_),
    .X(net303));
 sky130_fd_sc_hd__buf_8 fanout304 (.A(net305),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_16 fanout305 (.A(_1334_),
    .X(net305));
 sky130_fd_sc_hd__buf_8 fanout306 (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__buf_8 fanout307 (.A(_1317_),
    .X(net307));
 sky130_fd_sc_hd__buf_8 fanout308 (.A(_3494_),
    .X(net308));
 sky130_fd_sc_hd__buf_8 fanout309 (.A(_3494_),
    .X(net309));
 sky130_fd_sc_hd__buf_8 fanout310 (.A(_3418_),
    .X(net310));
 sky130_fd_sc_hd__buf_8 fanout311 (.A(_3418_),
    .X(net311));
 sky130_fd_sc_hd__buf_6 fanout312 (.A(_3417_),
    .X(net312));
 sky130_fd_sc_hd__buf_6 fanout313 (.A(_3417_),
    .X(net313));
 sky130_fd_sc_hd__buf_8 fanout314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_16 fanout315 (.A(net316),
    .X(net315));
 sky130_fd_sc_hd__buf_6 fanout317 (.A(_2732_),
    .X(net317));
 sky130_fd_sc_hd__buf_4 fanout318 (.A(_1702_),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_8 fanout319 (.A(_1690_),
    .X(net319));
 sky130_fd_sc_hd__buf_4 fanout320 (.A(_1679_),
    .X(net320));
 sky130_fd_sc_hd__buf_4 fanout321 (.A(_1667_),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_8 fanout322 (.A(_1655_),
    .X(net322));
 sky130_fd_sc_hd__buf_4 fanout323 (.A(_1644_),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_8 fanout324 (.A(_1633_),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_8 fanout325 (.A(_1624_),
    .X(net325));
 sky130_fd_sc_hd__buf_4 fanout326 (.A(_1596_),
    .X(net326));
 sky130_fd_sc_hd__buf_4 fanout327 (.A(_1584_),
    .X(net327));
 sky130_fd_sc_hd__buf_4 fanout328 (.A(_1575_),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_8 fanout329 (.A(_1564_),
    .X(net329));
 sky130_fd_sc_hd__buf_6 fanout330 (.A(_1548_),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_8 fanout331 (.A(_1535_),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_8 fanout332 (.A(_1523_),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_8 fanout333 (.A(_1510_),
    .X(net333));
 sky130_fd_sc_hd__buf_6 fanout334 (.A(_1498_),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_8 fanout335 (.A(_1487_),
    .X(net335));
 sky130_fd_sc_hd__buf_4 fanout336 (.A(_1475_),
    .X(net336));
 sky130_fd_sc_hd__buf_4 fanout337 (.A(_1463_),
    .X(net337));
 sky130_fd_sc_hd__buf_4 fanout338 (.A(_1452_),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_8 fanout339 (.A(_1442_),
    .X(net339));
 sky130_fd_sc_hd__buf_4 fanout340 (.A(_1432_),
    .X(net340));
 sky130_fd_sc_hd__buf_4 fanout341 (.A(_1420_),
    .X(net341));
 sky130_fd_sc_hd__buf_4 fanout342 (.A(_1407_),
    .X(net342));
 sky130_fd_sc_hd__buf_4 fanout343 (.A(_1396_),
    .X(net343));
 sky130_fd_sc_hd__buf_4 fanout344 (.A(_1366_),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_8 fanout345 (.A(_1355_),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_8 fanout346 (.A(_1343_),
    .X(net346));
 sky130_fd_sc_hd__buf_6 fanout347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__buf_6 fanout348 (.A(_1327_),
    .X(net348));
 sky130_fd_sc_hd__buf_6 fanout349 (.A(_1310_),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_4 fanout350 (.A(_1310_),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_8 fanout351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_8 fanout352 (.A(_1301_),
    .X(net352));
 sky130_fd_sc_hd__buf_12 fanout353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_16 fanout354 (.A(net355),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_8 fanout356 (.A(_2733_),
    .X(net356));
 sky130_fd_sc_hd__buf_4 fanout357 (.A(_2733_),
    .X(net357));
 sky130_fd_sc_hd__buf_8 fanout358 (.A(_2730_),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_8 fanout359 (.A(_2730_),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_8 fanout360 (.A(_2727_),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_8 fanout361 (.A(_2727_),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_8 fanout362 (.A(_2726_),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_8 fanout363 (.A(_2726_),
    .X(net363));
 sky130_fd_sc_hd__buf_6 fanout364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__buf_6 fanout365 (.A(_1323_),
    .X(net365));
 sky130_fd_sc_hd__buf_6 fanout366 (.A(net367),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_16 fanout367 (.A(_1341_),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_8 fanout368 (.A(_1316_),
    .X(net368));
 sky130_fd_sc_hd__buf_6 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_16 fanout370 (.A(_1315_),
    .X(net370));
 sky130_fd_sc_hd__buf_8 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__buf_12 fanout372 (.A(_1314_),
    .X(net372));
 sky130_fd_sc_hd__buf_8 fanout373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__buf_6 fanout374 (.A(_1284_),
    .X(net374));
 sky130_fd_sc_hd__buf_6 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__buf_8 fanout376 (.A(\U_DATAPATH.U_ID_EX.o_addr_src_EX ),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_16 fanout377 (.A(net2288),
    .X(net377));
 sky130_fd_sc_hd__buf_4 fanout378 (.A(net2288),
    .X(net378));
 sky130_fd_sc_hd__buf_8 fanout379 (.A(net2112),
    .X(net379));
 sky130_fd_sc_hd__buf_8 fanout380 (.A(net2112),
    .X(net380));
 sky130_fd_sc_hd__buf_8 fanout381 (.A(net2098),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_8 fanout382 (.A(net2098),
    .X(net382));
 sky130_fd_sc_hd__buf_8 fanout383 (.A(net2098),
    .X(net383));
 sky130_fd_sc_hd__buf_8 fanout384 (.A(net2098),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_4 fanout385 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_8 fanout386 (.A(net387),
    .X(net386));
 sky130_fd_sc_hd__buf_6 fanout387 (.A(net2096),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_8 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_8 fanout389 (.A(net2096),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_8 fanout390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_8 fanout391 (.A(net2096),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_8 fanout392 (.A(net395),
    .X(net392));
 sky130_fd_sc_hd__buf_2 fanout393 (.A(net395),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_8 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__buf_4 fanout395 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ),
    .X(net395));
 sky130_fd_sc_hd__buf_8 fanout396 (.A(net398),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_8 fanout397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__buf_4 fanout398 (.A(net400),
    .X(net398));
 sky130_fd_sc_hd__buf_8 fanout399 (.A(net400),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_8 fanout400 (.A(net2089),
    .X(net400));
 sky130_fd_sc_hd__buf_8 fanout401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__buf_8 fanout402 (.A(net406),
    .X(net402));
 sky130_fd_sc_hd__buf_8 fanout403 (.A(net406),
    .X(net403));
 sky130_fd_sc_hd__buf_8 fanout404 (.A(net406),
    .X(net404));
 sky130_fd_sc_hd__buf_4 fanout405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__buf_6 fanout406 (.A(net2297),
    .X(net406));
 sky130_fd_sc_hd__buf_8 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__buf_8 fanout408 (.A(net409),
    .X(net408));
 sky130_fd_sc_hd__buf_6 fanout409 (.A(net2286),
    .X(net409));
 sky130_fd_sc_hd__buf_8 fanout410 (.A(net414),
    .X(net410));
 sky130_fd_sc_hd__buf_8 fanout411 (.A(net414),
    .X(net411));
 sky130_fd_sc_hd__buf_8 fanout412 (.A(net414),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_8 fanout413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_16 fanout414 (.A(net2177),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_8 fanout415 (.A(net417),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_4 fanout416 (.A(net417),
    .X(net416));
 sky130_fd_sc_hd__buf_4 fanout417 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_8 fanout418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__buf_4 fanout419 (.A(net2174),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_8 fanout420 (.A(net421),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_8 fanout421 (.A(net2174),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_8 fanout422 (.A(net424),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_8 fanout423 (.A(net424),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_8 fanout424 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ),
    .X(net424));
 sky130_fd_sc_hd__buf_8 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__buf_8 fanout426 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net426));
 sky130_fd_sc_hd__buf_8 fanout427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__buf_4 fanout428 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net428));
 sky130_fd_sc_hd__buf_6 fanout429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__buf_8 fanout430 (.A(net434),
    .X(net430));
 sky130_fd_sc_hd__buf_8 fanout431 (.A(net434),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_4 fanout432 (.A(net434),
    .X(net432));
 sky130_fd_sc_hd__buf_8 fanout433 (.A(net434),
    .X(net433));
 sky130_fd_sc_hd__buf_8 fanout434 (.A(net2345),
    .X(net434));
 sky130_fd_sc_hd__buf_6 fanout435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__buf_6 fanout436 (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .X(net436));
 sky130_fd_sc_hd__buf_4 fanout437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__buf_4 fanout438 (.A(_0069_),
    .X(net438));
 sky130_fd_sc_hd__buf_4 fanout439 (.A(_0069_),
    .X(net439));
 sky130_fd_sc_hd__buf_2 fanout440 (.A(_0069_),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_4 fanout441 (.A(_0069_),
    .X(net441));
 sky130_fd_sc_hd__buf_2 fanout442 (.A(_0069_),
    .X(net442));
 sky130_fd_sc_hd__buf_4 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__buf_4 fanout444 (.A(net448),
    .X(net444));
 sky130_fd_sc_hd__buf_4 fanout445 (.A(net448),
    .X(net445));
 sky130_fd_sc_hd__buf_4 fanout446 (.A(net448),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_8 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_4 fanout448 (.A(_0069_),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_4 fanout449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__buf_4 fanout450 (.A(net463),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_4 fanout451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__buf_4 fanout452 (.A(net463),
    .X(net452));
 sky130_fd_sc_hd__buf_4 fanout453 (.A(net463),
    .X(net453));
 sky130_fd_sc_hd__buf_4 fanout454 (.A(net463),
    .X(net454));
 sky130_fd_sc_hd__buf_4 fanout455 (.A(net463),
    .X(net455));
 sky130_fd_sc_hd__buf_4 fanout456 (.A(net463),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_4 fanout457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__buf_4 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_8 fanout459 (.A(net463),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_8 fanout460 (.A(net462),
    .X(net460));
 sky130_fd_sc_hd__buf_4 fanout461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__buf_4 fanout462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__buf_6 fanout463 (.A(_0069_),
    .X(net463));
 sky130_fd_sc_hd__buf_8 fanout464 (.A(net466),
    .X(net464));
 sky130_fd_sc_hd__buf_4 fanout465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__buf_6 fanout466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__buf_8 fanout467 (.A(net63),
    .X(net467));
 sky130_fd_sc_hd__buf_8 fanout468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__buf_8 fanout469 (.A(net63),
    .X(net469));
 sky130_fd_sc_hd__buf_8 fanout470 (.A(net63),
    .X(net470));
 sky130_fd_sc_hd__buf_8 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__buf_4 fanout472 (.A(net63),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[8] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0550_),
    .X(net553));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold100 (.A(_0853_),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(_0481_),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(_1161_),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(_0340_),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(_1062_),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(_0482_),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[13] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(_1214_),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(_0386_),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(_0895_),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(_0360_),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(_1012_),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0836_),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(_1207_),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(_1177_),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(_0975_),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(_0979_),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(_0490_),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[19] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(_0327_),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(_1073_),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(_1000_),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(_0500_),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(_0374_),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_0302_),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(_0394_),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(_0448_),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(_0966_),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(_0976_),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(_1213_),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[27] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(_0999_),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(_1236_),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(_0337_),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(_1221_),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(_1238_),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0567_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(_1171_),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(_0411_),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(_1239_),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(_1223_),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(_0505_),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[25] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(_0344_),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(_0405_),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(_1197_),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(_0424_),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(_0390_),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0710_),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(_1033_),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(_0498_),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(_1072_),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(_1147_),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(_1230_),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[11] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(_0496_),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(_0486_),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(_1148_),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(_0362_),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(_0501_),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[2] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0802_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(_1225_),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(_0503_),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(_1194_),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(_1104_),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(_0399_),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[20] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(_0488_),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(_0383_),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(_1178_),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(_1163_),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(_0412_),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0811_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(_1034_),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(_1182_),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(_1153_),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(_0436_),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(_0476_),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[27] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(_0328_),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(_0473_),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(_1219_),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(_0964_),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(_0402_),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_0712_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(_1228_),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(_1020_),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(_0404_),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(_1075_),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(_0493_),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[29] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(_0358_),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(_0492_),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(_1160_),
    .X(net1697));
 sky130_fd_sc_hd__clkbuf_8 hold1155 (.A(net2205),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(_3612_),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(_1264_),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(_0985_),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_0539_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(_1155_),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(_1049_),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(_1224_),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(_1027_),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(_1170_),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(net116),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(_0329_),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(_1184_),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(_0470_),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(_1231_),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_0685_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(_0897_),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(_0318_),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(_0913_),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(_0475_),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(_0941_),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[16] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(_1243_),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(_1037_),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(_0345_),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(_1183_),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(_1146_),
    .X(net1741));
 sky130_fd_sc_hd__clkbuf_2 hold1199 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[28] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0542_),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0807_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(_1268_),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(_1150_),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(_0935_),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(_1165_),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(_0914_),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[14] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(_0980_),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(_1179_),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(_1007_),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(_1154_),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(_1157_),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0837_),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(_1023_),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(_1045_),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(_1195_),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(_0953_),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(_1151_),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[3] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(_1028_),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(_0444_),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(_1039_),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(_1164_),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(net102),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(_0946_),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0688_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(_1167_),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(_0951_),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(_1201_),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(_1185_),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(_1172_),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[15] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(_1169_),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(_1048_),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(net109),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(_0922_),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(_0926_),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_0838_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(_0923_),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(_0489_),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(_1196_),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(_1051_),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(_1168_),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ),
    .X(net1812));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold127 (.A(net2357),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(_0937_),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(_0504_),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(_1200_),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(_1019_),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(_1036_),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\U_DATAPATH.U_EX_MEM.o_result_src_M[1] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(_1173_),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(_0925_),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(_0408_),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(_1162_),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(_0929_),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0194_),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(_1189_),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(_0942_),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(_1158_),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(_0936_),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(_0928_),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[20] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[9] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(_1186_),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(_1191_),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(_0943_),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(_1159_),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(net118),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(_0940_),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_0832_),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(_1204_),
    .X(net1854));
 sky130_fd_sc_hd__buf_1 hold1312 (.A(net2359),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(_1174_),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(_1029_),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(_1031_),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[5] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(_1199_),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(_1206_),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(_0939_),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(_0684_),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(_1024_),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_0828_),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(_1190_),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[21] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(_0244_),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(_0933_),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[0] ),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(_2683_),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(_0651_),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(_1192_),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[14] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(_1038_),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(_1152_),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[30] ),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(_0253_),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(_1046_),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(_0938_),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0699_),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(_0927_),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(_0945_),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(_0950_),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(_1025_),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(net105),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[10] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(_1035_),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(_1205_),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(_0952_),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(_0949_),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(_0947_),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0695_),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(_1044_),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(_1043_),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(_0930_),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(_1193_),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(_1156_),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[22] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(_1041_),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(_1042_),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(_1030_),
    .X(net1927));
 sky130_fd_sc_hd__clkbuf_2 hold1385 (.A(net2084),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(_0948_),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(_1018_),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_0813_),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(_0478_),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(_1198_),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(_0931_),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(_1166_),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(_0932_),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0705_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[26] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(net108),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(net107),
    .X(net1944));
 sky130_fd_sc_hd__clkbuf_4 hold1402 (.A(net2368),
    .X(net1945));
 sky130_fd_sc_hd__clkbuf_4 hold1403 (.A(_3605_),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(_1258_),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(_1026_),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(_0934_),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_0817_),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(_1144_),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[28] ),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(_0251_),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(_1032_),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(_1187_),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(net119),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(_1202_),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[17] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(_0944_),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(_1040_),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(_1083_),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(_1188_),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[13] ),
    .X(net1971));
 sky130_fd_sc_hd__buf_2 hold1429 (.A(net2358),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_0840_),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(_3597_),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(_1250_),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(_1180_),
    .X(net1976));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1434 (.A(net73),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(_1047_),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(_1022_),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[11] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(_0791_),
    .X(net1983));
 sky130_fd_sc_hd__buf_2 hold1441 (.A(net2365),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(_0792_),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(\U_DATAPATH.U_EX_MEM.i_result_src_EX[0] ),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[22] ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[14] ),
    .X(net1989));
 sky130_fd_sc_hd__clkbuf_8 hold1447 (.A(net2215),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(_3610_),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[6] ),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_0834_),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[5] ),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(_1117_),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(net123),
    .X(net1995));
 sky130_fd_sc_hd__clkbuf_2 hold1453 (.A(net2363),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(net114),
    .X(net1997));
 sky130_fd_sc_hd__clkbuf_8 hold1455 (.A(net2197),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(_3611_),
    .X(net1999));
 sky130_fd_sc_hd__buf_1 hold1457 (.A(net2369),
    .X(net2000));
 sky130_fd_sc_hd__clkbuf_8 hold1458 (.A(net2125),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(_3595_),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[6] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(_1248_),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[3] ),
    .X(net2004));
 sky130_fd_sc_hd__buf_1 hold1462 (.A(net2374),
    .X(net2005));
 sky130_fd_sc_hd__clkbuf_2 hold1463 (.A(net2372),
    .X(net2006));
 sky130_fd_sc_hd__buf_1 hold1464 (.A(net2370),
    .X(net2007));
 sky130_fd_sc_hd__clkbuf_2 hold1465 (.A(net2371),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(_0683_),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(net101),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(net121),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0797_),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[9] ),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(_1121_),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[15] ),
    .X(net2015));
 sky130_fd_sc_hd__buf_1 hold1473 (.A(net2373),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[7] ),
    .X(net2017));
 sky130_fd_sc_hd__clkbuf_2 hold1475 (.A(net2361),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(_3598_),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(_1251_),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[23] ),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(_1135_),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[24] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[16] ),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[19] ),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(_1949_),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(_1960_),
    .X(net2026));
 sky130_fd_sc_hd__buf_1 hold1484 (.A(net2376),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(_1895_),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[27] ),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[0] ),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[29] ),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(_2040_),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_0709_),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(net66),
    .X(net2033));
 sky130_fd_sc_hd__buf_2 hold1491 (.A(net2360),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(net126),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[31] ),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(\U_DATAPATH.U_EX_MEM.i_mem_write_EX ),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(_0790_),
    .X(net2039));
 sky130_fd_sc_hd__buf_1 hold1497 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[28] ),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(_2026_),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(_2038_),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[22] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[19] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(_2039_),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[10] ),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(_1122_),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(net104),
    .X(net2046));
 sky130_fd_sc_hd__clkbuf_2 hold1504 (.A(net2364),
    .X(net2047));
 sky130_fd_sc_hd__clkbuf_2 hold1505 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(_2679_),
    .X(net2049));
 sky130_fd_sc_hd__clkbuf_2 hold1507 (.A(_2680_),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(_3609_),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[26] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_0842_),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(_2013_),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[4] ),
    .X(net2054));
 sky130_fd_sc_hd__buf_1 hold1512 (.A(net2362),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(_2004_),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(_2005_),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(net65),
    .X(net2058));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1516 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[24] ),
    .X(net2059));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1517 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[11] ),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[8] ),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[16] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(_0789_),
    .X(net2063));
 sky130_fd_sc_hd__buf_1 hold1521 (.A(net2367),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(_1132_),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(net75),
    .X(net2066));
 sky130_fd_sc_hd__clkbuf_2 hold1524 (.A(net2377),
    .X(net2067));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1525 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[17] ),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(net129),
    .X(net2069));
 sky130_fd_sc_hd__clkbuf_2 hold1527 (.A(net2380),
    .X(net2070));
 sky130_fd_sc_hd__clkbuf_2 hold1528 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .X(net2071));
 sky130_fd_sc_hd__clkbuf_4 hold1529 (.A(_2135_),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_0701_),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_4 hold1530 (.A(net2389),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .X(net2074));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1532 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(_1917_),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(_1928_),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(_1929_),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(_1931_),
    .X(net2079));
 sky130_fd_sc_hd__buf_1 hold1537 (.A(net2375),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(_1176_),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[18] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(\U_CONTROL_UNIT.i_jump_EX ),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(net90),
    .X(net2084));
 sky130_fd_sc_hd__clkbuf_8 hold1542 (.A(net174),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(_1145_),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(net100),
    .X(net2088));
 sky130_fd_sc_hd__buf_1 hold1546 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(_3603_),
    .X(net2090));
 sky130_fd_sc_hd__buf_4 hold1548 (.A(net2384),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(_3593_),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_0703_),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(_0924_),
    .X(net2094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(net111),
    .X(net2095));
 sky130_fd_sc_hd__buf_2 hold1553 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(_3602_),
    .X(net2097));
 sky130_fd_sc_hd__clkbuf_4 hold1555 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(_3601_),
    .X(net2099));
 sky130_fd_sc_hd__buf_1 hold1557 (.A(net2388),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(_0225_),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ),
    .X(net2102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[25] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(_1021_),
    .X(net2103));
 sky130_fd_sc_hd__clkbuf_2 hold1561 (.A(net2378),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(\U_DATAPATH.U_EX_MEM.i_funct3_EX[2] ),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(net122),
    .X(net2106));
 sky130_fd_sc_hd__buf_2 hold1564 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[3] ),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(_0647_),
    .X(net2108));
 sky130_fd_sc_hd__buf_1 hold1566 (.A(net2366),
    .X(net2109));
 sky130_fd_sc_hd__clkbuf_4 hold1567 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[24] ),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(_3599_),
    .X(net2111));
 sky130_fd_sc_hd__buf_2 hold1569 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .X(net2112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_0816_),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(_3600_),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(_1181_),
    .X(net2115));
 sky130_fd_sc_hd__clkbuf_2 hold1573 (.A(net2381),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(net125),
    .X(net2117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(net120),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(net112),
    .X(net2119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(net124),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(\U_CONTROL_UNIT.i_branch_EX ),
    .X(net2121));
 sky130_fd_sc_hd__clkbuf_2 hold1579 (.A(net183),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[23] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(net106),
    .X(net2123));
 sky130_fd_sc_hd__clkbuf_2 hold1581 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(_2134_),
    .X(net2125));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1583 (.A(net2391),
    .X(net2126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(_1149_),
    .X(net2128));
 sky130_fd_sc_hd__buf_1 hold1586 (.A(net2390),
    .X(net2129));
 sky130_fd_sc_hd__clkbuf_2 hold1587 (.A(net2382),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[11] ),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ),
    .X(net2132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_0814_),
    .X(net702));
 sky130_fd_sc_hd__buf_1 hold1590 (.A(_1944_),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(_1956_),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(_1957_),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[1] ),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(_1788_),
    .X(net2137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(_1789_),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(_0652_),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[25] ),
    .X(net2140));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1598 (.A(_1476_),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(net115),
    .X(net2142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0845_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[3] ),
    .X(net703));
 sky130_fd_sc_hd__buf_1 hold1600 (.A(net2383),
    .X(net2143));
 sky130_fd_sc_hd__clkbuf_4 hold1601 (.A(net2386),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[12] ),
    .X(net2145));
 sky130_fd_sc_hd__buf_1 hold1603 (.A(_1691_),
    .X(net2146));
 sky130_fd_sc_hd__buf_1 hold1604 (.A(net2387),
    .X(net2147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[18] ),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(_1935_),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(_1947_),
    .X(net2150));
 sky130_fd_sc_hd__clkbuf_2 hold1608 (.A(net2379),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(net91),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_0826_),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_4 hold1610 (.A(net2385),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(_1782_),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(_1784_),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(_1798_),
    .X(net2157));
 sky130_fd_sc_hd__clkbuf_2 hold1615 (.A(net88),
    .X(net2158));
 sky130_fd_sc_hd__clkbuf_4 hold1616 (.A(net80),
    .X(net2159));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1617 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(_1835_),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(_1847_),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[19] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(_1848_),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(_1881_),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(_1892_),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(_1893_),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(net74),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ),
    .X(net2169));
 sky130_fd_sc_hd__clkbuf_2 hold1627 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(_1816_),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(_1828_),
    .X(net2172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_0810_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(_1829_),
    .X(net2173));
 sky130_fd_sc_hd__clkbuf_2 hold1631 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(_1825_),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ),
    .X(net2177));
 sky130_fd_sc_hd__buf_2 hold1635 (.A(net83),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(net117),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[31] ),
    .X(net2180));
 sky130_fd_sc_hd__buf_1 hold1638 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(_1972_),
    .X(net2182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[9] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(_1984_),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(_1985_),
    .X(net2184));
 sky130_fd_sc_hd__clkbuf_2 hold1642 (.A(net78),
    .X(net2185));
 sky130_fd_sc_hd__buf_1 hold1643 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(_2017_),
    .X(net2187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(_2029_),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[10] ),
    .X(net2189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(_1863_),
    .X(net2190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(_1875_),
    .X(net2191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(_1876_),
    .X(net2192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_0694_),
    .X(net708));
 sky130_fd_sc_hd__buf_1 hold1650 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(_1898_),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(_1911_),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(_1912_),
    .X(net2196));
 sky130_fd_sc_hd__buf_2 hold1654 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .X(net2197));
 sky130_fd_sc_hd__clkbuf_2 hold1655 (.A(net85),
    .X(net2198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1656 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(_1925_),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .X(net2202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[8] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[21] ),
    .X(net2203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[19] ),
    .X(net2204));
 sky130_fd_sc_hd__clkbuf_2 hold1662 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ),
    .X(net2205));
 sky130_fd_sc_hd__buf_1 hold1663 (.A(_3570_),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(_1209_),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[26] ),
    .X(net2208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[5] ),
    .X(net2209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ),
    .X(net2210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(_1981_),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(_1993_),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_0799_),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(_1994_),
    .X(net2213));
 sky130_fd_sc_hd__buf_1 hold1671 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(_2035_),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(_2045_),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(_2046_),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[29] ),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(net86),
    .X(net2221));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1679 (.A(_1368_),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[3] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[10] ),
    .X(net2223));
 sky130_fd_sc_hd__clkbuf_2 hold1681 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(_1844_),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1684 (.A(_1908_),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(_1920_),
    .X(net2228));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1686 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(_1811_),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1688 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .X(net2231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(net183),
    .X(net2232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_0286_),
    .X(net712));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1690 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ),
    .X(net2233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(_2008_),
    .X(net2234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(_2020_),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[0] ),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[13] ),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(_1887_),
    .X(net2238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(_1901_),
    .X(net2239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ),
    .X(net2240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(_1854_),
    .X(net2241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(net128),
    .X(net2242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[28] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[8] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ),
    .X(net2243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(_1953_),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(_1966_),
    .X(net2245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(_1967_),
    .X(net2246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[31] ),
    .X(net2247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(_2051_),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(_2052_),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[7] ),
    .X(net2250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(_1577_),
    .X(net2251));
 sky130_fd_sc_hd__buf_1 hold1709 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[3] ),
    .X(net2252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_0693_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[17] ),
    .X(net2253));
 sky130_fd_sc_hd__buf_1 hold1711 (.A(_0769_),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[14] ),
    .X(net2255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[8] ),
    .X(net2256));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1714 (.A(_1645_),
    .X(net2257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[4] ),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1716 (.A(_1805_),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[29] ),
    .X(net2260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(_3379_),
    .X(net2261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(_0746_),
    .X(net2262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[21] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1720 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(_1963_),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(_1975_),
    .X(net2265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[23] ),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[6] ),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[13] ),
    .X(net2269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1727 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[28] ),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(_1351_),
    .X(net2271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1729 (.A(_0745_),
    .X(net2272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_0706_),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[20] ),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[28] ),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1732 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[27] ),
    .X(net2275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[11] ),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(_3411_),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[15] ),
    .X(net2279));
 sky130_fd_sc_hd__buf_1 hold1737 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[16] ),
    .X(net2280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ),
    .X(net2281));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1739 (.A(_1478_),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[22] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(_1479_),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(_3313_),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(_0742_),
    .X(net2285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .X(net2286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1744 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .X(net2287));
 sky130_fd_sc_hd__clkbuf_2 hold1745 (.A(\U_DATAPATH.U_ID_EX.o_alu_src_EX ),
    .X(net2288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1746 (.A(_1698_),
    .X(net2289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1747 (.A(_0729_),
    .X(net2290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1748 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[24] ),
    .X(net2291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[18] ),
    .X(net2292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_0707_),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1750 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(_1447_),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(_1448_),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1753 (.A(_0739_),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ),
    .X(net2297));
 sky130_fd_sc_hd__buf_1 hold1755 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[2] ),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1756 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[4] ),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ),
    .X(net2300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ),
    .X(net2301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1759 (.A(_1506_),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[23] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1760 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ),
    .X(net2303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1761 (.A(_0733_),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1762 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1763 (.A(_0734_),
    .X(net2306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1764 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[23] ),
    .X(net2307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1765 (.A(_0740_),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1766 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .X(net2309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1767 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[21] ),
    .X(net2310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1768 (.A(_0738_),
    .X(net2311));
 sky130_fd_sc_hd__buf_1 hold1769 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[30] ),
    .X(net2312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_0846_),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1770 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1771 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ),
    .X(net2314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1772 (.A(_0730_),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1773 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[22] ),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1774 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[19] ),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1775 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[25] ),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1776 (.A(_1997_),
    .X(net2319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1777 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[7] ),
    .X(net2320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1778 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[14] ),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1779 (.A(_0731_),
    .X(net2322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[7] ),
    .X(net721));
 sky130_fd_sc_hd__buf_1 hold1780 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1781 (.A(_1771_),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1782 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[2] ),
    .X(net2325));
 sky130_fd_sc_hd__clkbuf_2 hold1783 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ),
    .X(net2326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1784 (.A(_1774_),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1785 (.A(_2740_),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1786 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ),
    .X(net2329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1787 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[27] ),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1788 (.A(_1516_),
    .X(net2331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1789 (.A(_0744_),
    .X(net2332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_0830_),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1790 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[20] ),
    .X(net2333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1791 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[24] ),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1792 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[1] ),
    .X(net2335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1793 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ),
    .X(net2336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1794 (.A(_3018_),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1795 (.A(_0726_),
    .X(net2338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1796 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[8] ),
    .X(net2339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1797 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[5] ),
    .X(net2340));
 sky130_fd_sc_hd__buf_1 hold1798 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1799 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[26] ),
    .X(net2342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0851_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[24] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1800 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[15] ),
    .X(net2343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1801 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[9] ),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1802 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net2345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1803 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[10] ),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1804 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[18] ),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1805 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[11] ),
    .X(net2348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1806 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[4] ),
    .X(net2349));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1807 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ),
    .X(net2350));
 sky130_fd_sc_hd__buf_1 hold1808 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[3] ),
    .X(net2351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1809 (.A(net110),
    .X(net2352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_0815_),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1810 (.A(net103),
    .X(net2353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1811 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ),
    .X(net2354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1812 (.A(net113),
    .X(net2355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1813 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .X(net2356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1814 (.A(net87),
    .X(net2357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1815 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[26] ),
    .X(net2358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1816 (.A(net68),
    .X(net2359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1817 (.A(net93),
    .X(net2360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1818 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[25] ),
    .X(net2361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1819 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[25] ),
    .X(net2362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[5] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1820 (.A(net84),
    .X(net2363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1821 (.A(net71),
    .X(net2364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1822 (.A(net89),
    .X(net2365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1823 (.A(\U_DATAPATH.U_EX_MEM.o_reg_write_M ),
    .X(net2366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1824 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[20] ),
    .X(net2367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1825 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[31] ),
    .X(net2368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1826 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ),
    .X(net2369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1827 (.A(net64),
    .X(net2370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1828 (.A(net94),
    .X(net2371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1829 (.A(net81),
    .X(net2372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_0545_),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1830 (.A(net79),
    .X(net2373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1831 (.A(net77),
    .X(net2374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1832 (.A(net76),
    .X(net2375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1833 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[12] ),
    .X(net2376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1834 (.A(net92),
    .X(net2377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1835 (.A(net95),
    .X(net2378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1836 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[1] ),
    .X(net2379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1837 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[18] ),
    .X(net2380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1838 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[27] ),
    .X(net2381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1839 (.A(net67),
    .X(net2382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[17] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1840 (.A(net82),
    .X(net2383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1841 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ),
    .X(net2384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1842 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[2] ),
    .X(net2385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1843 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ),
    .X(net2386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1844 (.A(net69),
    .X(net2387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1845 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[2] ),
    .X(net2388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1846 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[29] ),
    .X(net2389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1847 (.A(net70),
    .X(net2390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1848 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[19] ),
    .X(net2391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_0808_),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[17] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_0702_),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[12] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_0697_),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[20] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[7] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_0798_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[31] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_0716_),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[28] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_0713_),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\U_DATAPATH.U_EX_MEM.i_reg_write_EX ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_0751_),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[8] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_0548_),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0291_),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0843_),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_0686_),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(net2118),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[2] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_0825_),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\U_DATAPATH.U_EX_MEM.i_funct3_EX[1] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_0786_),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[12] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_0803_),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[23] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[18] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0708_),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[29] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_0714_),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[30] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_0715_),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[18] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_0841_),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[24] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_0307_),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[8] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0809_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_0518_),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[26] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_0536_),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[30] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_0821_),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[28] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_0819_),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[2] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_0793_),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[31] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[19] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_0541_),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[25] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0535_),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[23] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_0306_),
    .X(net777));
 sky130_fd_sc_hd__buf_1 hold235 (.A(net2033),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(net2352),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[11] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_0696_),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[13] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0704_),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0296_),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_1050_),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_1084_),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[9] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_0549_),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_0477_),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[15] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[0] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_0555_),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_0956_),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(net2142),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_1052_),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[19] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_0529_),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_0413_),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0823_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[27] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_0537_),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_0954_),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[13] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(_0523_),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(net2353),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_0890_),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[31] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_0382_),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[30] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_0570_),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[16] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_0299_),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[31] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_0314_),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[24] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_0534_),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[11] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0854_),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_0551_),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[7] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_0290_),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[12] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_0295_),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[27] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_0310_),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[14] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_0297_),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[11] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[10] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_0521_),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[12] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_0522_),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[30] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_0313_),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[4] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_0514_),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[7] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_0547_),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[6] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[2] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0833_),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_0546_),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[11] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_0294_),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[28] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_0311_),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[20] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_0560_),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[6] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_0289_),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[15] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_0443_),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[22] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_0305_),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[15] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_0525_),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[18] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_0301_),
    .X(net859));
 sky130_fd_sc_hd__buf_2 hold317 (.A(net2221),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[21] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(_0304_),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0806_),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[31] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(_0571_),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[5] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(_0288_),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(_0989_),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_0350_),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[21] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_0531_),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[13] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_0891_),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[28] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_0568_),
    .X(net876));
 sky130_fd_sc_hd__buf_2 hold334 (.A(net2030),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[13] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_0553_),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[4] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_0287_),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0698_),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_0516_),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[14] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_0554_),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[5] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_0515_),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[20] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_0303_),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[15] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_0298_),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[27] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_0921_),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[3] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_0513_),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[26] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_0309_),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(net72),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(_0917_),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[10] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(_0520_),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0850_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(_0379_),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(_0907_),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(_1067_),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[23] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(_0563_),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(_0986_),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[12] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(_0414_),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[23] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(_0533_),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(_1106_),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[9] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(_0519_),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[2] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(_0285_),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0552_),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(_0455_),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(_0366_),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(_1005_),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(net2355),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[7] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_0517_),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[4] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_1113_),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_0391_),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(_0315_),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_0409_),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_1082_),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0687_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0689_),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_1078_),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_1109_),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[25] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_0308_),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[22] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_0532_),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_0451_),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[5] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_0439_),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_0446_),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[25] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_0565_),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[9] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_0292_),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[24] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_0564_),
    .X(net961));
 sky130_fd_sc_hd__buf_1 hold419 (.A(net2058),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0796_),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(_1066_),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(_0346_),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(_0364_),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[4] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(_0544_),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[17] ),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(_0300_),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[3] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(_1074_),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[10] ),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(_0293_),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(_0892_),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(_0978_),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(_0982_),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0794_),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[28] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(_0538_),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(_1081_),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(_0899_),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(_0377_),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(_1110_),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[5] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(_1069_),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(_0317_),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(_0396_),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(_0427_),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(_0460_),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0690_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(_0415_),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(_1016_),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(_0973_),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(_0992_),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\U_DATAPATH.U_IF_ID.i_pc_IF[29] ),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(_0312_),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[29] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(_0423_),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(_0352_),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[22] ),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(_0562_),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(_0965_),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(_0389_),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0852_),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_0375_),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(_0316_),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(_1101_),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[16] ),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(_0526_),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[18] ),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(_0528_),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[27] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(_0384_),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(_0969_),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(_0400_),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(_0371_),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[14] ),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(_0524_),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[16] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0818_),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(_0433_),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(_1013_),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(_0348_),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(_0458_),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(_0900_),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[31] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(_1240_),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(_0369_),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(_0355_),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(_0403_),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[21] ),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(_0561_),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0822_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(_0464_),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[29] ),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(_0569_),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(_0909_),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(_0479_),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(_0957_),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\U_DATAPATH.U_EX_MEM.i_funct3_EX[0] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(_0319_),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(_0959_),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[18] ),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(_0558_),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(_1064_),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(_1102_),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0785_),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(_0474_),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[26] ),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(_0566_),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(_1234_),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(_1055_),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(_1108_),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[9] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(_0343_),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[19] ),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(_0559_),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(_0445_),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(_0332_),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(_0351_),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0800_),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(_1217_),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(_0428_),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(_0372_),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(_1095_),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(_0419_),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[6] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(_0323_),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(_0321_),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[2] ),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(_0512_),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(_0334_),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(_0984_),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0691_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(_0901_),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[20] ),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(_0530_),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(_0967_),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(_0341_),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(_0420_),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[7] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(_0336_),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[3] ),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(_0543_),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(_1103_),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(_0898_),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(_1094_),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0556_),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0692_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(_1098_),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(_0908_),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(_0893_),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(_0903_),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(_0370_),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[13] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(_1215_),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(_0447_),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(_1059_),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(_0426_),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(_1014_),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0804_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(_1105_),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(_0325_),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(_0338_),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(_0357_),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(_0494_),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[12] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(_0963_),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(_0422_),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(_0440_),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(_0378_),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(_0906_),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0835_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(_0918_),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(_0997_),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(_0962_),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(_0915_),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(_1017_),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[17] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(_0376_),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(_0454_),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(_0896_),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(_0988_),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(_0381_),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0527_),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(_0960_),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(_0994_),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(_0974_),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(_1220_),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(_1015_),
    .X(net1212));
 sky130_fd_sc_hd__buf_1 hold67 (.A(\U_DATAPATH.U_EX_MEM.i_result_src_EX[1] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(_0904_),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(_0330_),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(_0380_),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(_0385_),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(_0971_),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0750_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(_0459_),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(_1099_),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[17] ),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(_0557_),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(_0483_),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(_0359_),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[8] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(_0485_),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(_0353_),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(_0995_),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(_0356_),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(_1065_),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[1] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0831_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(_1089_),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(_0911_),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(_0453_),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(_0502_),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(_0919_),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[15] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(_0471_),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(_0491_),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(_0450_),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(_1056_),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(_0418_),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0700_),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(_0387_),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(_1227_),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(_0397_),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(_1079_),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(_1107_),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[6] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(_1008_),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(_0894_),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(_1004_),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(_0438_),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[30] ),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(_0540_),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0829_),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(_0430_),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(_0410_),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(_0395_),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(_1216_),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(_0442_),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[14] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(_0905_),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(_0987_),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(_1093_),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(_0468_),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(_1097_),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0805_),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(_0406_),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(_1086_),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(_0466_),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(_0977_),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(_1096_),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[25] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(_0910_),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(_1085_),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(_0361_),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(_0435_),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(_0902_),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0848_),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(_0449_),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(_0499_),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(_0425_),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(_0506_),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(_1112_),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[4] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(_1071_),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(_0991_),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(_0452_),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(_0920_),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(_1232_),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0824_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0827_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(_1010_),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(_0421_),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(_0368_),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(_0484_),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(_0333_),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[10] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(_0373_),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(_0457_),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(_0363_),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(_1090_),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(_0367_),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0801_),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(_1088_),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(_0388_),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(_0432_),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(_0407_),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(_0968_),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[4] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(_0441_),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(_1063_),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(_1226_),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(_1237_),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(_0349_),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0795_),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(_0996_),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(_1001_),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(_1054_),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(_1087_),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(_0469_),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[21] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(_0998_),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(_0480_),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(_1011_),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(_0429_),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(_1111_),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0812_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(_1218_),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(_0993_),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(_0463_),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(_0461_),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(_0434_),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[16] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(_0912_),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(_1003_),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(net127),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(_0467_),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(_1241_),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0839_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(_1070_),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(_0393_),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(_1222_),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(_1058_),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(_0326_),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[21] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(_0487_),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(_1077_),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(_0990_),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(_1002_),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(_0398_),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[10] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0844_),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(_1203_),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(_0961_),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(_0354_),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(_0472_),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(_1235_),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\U_DATAPATH.U_EX_MEM.o_result_src_M[0] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(_1060_),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(_0981_),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(_0955_),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(_0324_),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(_1009_),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0193_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(_0322_),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(_0342_),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(_0431_),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(_0495_),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(_1053_),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[26] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(_1233_),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(_0462_),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[29] ),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(_0820_),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(_0417_),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(_0331_),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0711_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(_1229_),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(_0972_),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(_1091_),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(_0320_),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(_0983_),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[26] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(_1068_),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(_0465_),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(_0339_),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(_0970_),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(_0392_),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0849_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(_0416_),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(_0958_),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(_0365_),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(_1061_),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(_0401_),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[24] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(_1244_),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(_1080_),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(_0335_),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(_0456_),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(_0347_),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0847_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(_0916_),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(_1092_),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(_0437_),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(_1175_),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(_1100_),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[30] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(_1057_),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(_0497_),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(_1076_),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(_1242_),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(_1006_),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ),
    .X(net1542));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(i_instr_ID[10]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(i_instr_ID[19]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(i_instr_ID[20]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(i_instr_ID[21]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(i_instr_ID[22]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(i_instr_ID[23]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(i_instr_ID[24]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(i_instr_ID[25]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(i_instr_ID[26]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(i_instr_ID[27]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(i_instr_ID[28]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(i_instr_ID[11]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(i_instr_ID[29]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(i_instr_ID[2]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(i_instr_ID[30]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(i_instr_ID[31]),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input24 (.A(i_instr_ID[3]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(i_instr_ID[4]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(i_instr_ID[5]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(i_instr_ID[6]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(i_instr_ID[7]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(i_instr_ID[8]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(i_instr_ID[12]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(i_instr_ID[9]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(i_read_data_M[0]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(i_read_data_M[10]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(i_read_data_M[11]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(i_read_data_M[12]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input35 (.A(i_read_data_M[13]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(i_read_data_M[14]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input37 (.A(i_read_data_M[15]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(i_read_data_M[16]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 input39 (.A(i_read_data_M[17]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input4 (.A(i_instr_ID[13]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(i_read_data_M[18]),
    .X(net40));
 sky130_fd_sc_hd__buf_2 input41 (.A(i_read_data_M[19]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(i_read_data_M[1]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 input43 (.A(i_read_data_M[20]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(i_read_data_M[21]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(i_read_data_M[22]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(i_read_data_M[23]),
    .X(net46));
 sky130_fd_sc_hd__buf_4 input47 (.A(i_read_data_M[24]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(i_read_data_M[25]),
    .X(net48));
 sky130_fd_sc_hd__buf_4 input49 (.A(i_read_data_M[26]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input5 (.A(i_instr_ID[14]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input50 (.A(i_read_data_M[27]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(i_read_data_M[28]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(i_read_data_M[29]),
    .X(net52));
 sky130_fd_sc_hd__buf_4 input53 (.A(i_read_data_M[2]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(i_read_data_M[30]),
    .X(net54));
 sky130_fd_sc_hd__dlymetal6s2s_1 input55 (.A(i_read_data_M[31]),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(i_read_data_M[3]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(i_read_data_M[4]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(i_read_data_M[5]),
    .X(net58));
 sky130_fd_sc_hd__buf_2 input59 (.A(i_read_data_M[6]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(i_instr_ID[15]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(i_read_data_M[7]),
    .X(net60));
 sky130_fd_sc_hd__dlymetal6s2s_1 input61 (.A(i_read_data_M[8]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(i_read_data_M[9]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_8 input63 (.A(rst),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input7 (.A(i_instr_ID[16]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(i_instr_ID[17]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(i_instr_ID[18]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 max_cap316 (.A(_3412_),
    .X(net316));
 sky130_fd_sc_hd__buf_4 max_cap355 (.A(_1300_),
    .X(net355));
 sky130_fd_sc_hd__buf_12 output100 (.A(net100),
    .X(o_pc_IF[10]));
 sky130_fd_sc_hd__buf_12 output101 (.A(net101),
    .X(o_pc_IF[11]));
 sky130_fd_sc_hd__buf_12 output102 (.A(net102),
    .X(o_pc_IF[12]));
 sky130_fd_sc_hd__buf_12 output103 (.A(net103),
    .X(o_pc_IF[13]));
 sky130_fd_sc_hd__buf_12 output104 (.A(net104),
    .X(o_pc_IF[14]));
 sky130_fd_sc_hd__buf_12 output105 (.A(net105),
    .X(o_pc_IF[15]));
 sky130_fd_sc_hd__buf_12 output106 (.A(net106),
    .X(o_pc_IF[16]));
 sky130_fd_sc_hd__buf_12 output107 (.A(net107),
    .X(o_pc_IF[17]));
 sky130_fd_sc_hd__buf_12 output108 (.A(net108),
    .X(o_pc_IF[18]));
 sky130_fd_sc_hd__buf_12 output109 (.A(net109),
    .X(o_pc_IF[19]));
 sky130_fd_sc_hd__buf_12 output110 (.A(net110),
    .X(o_pc_IF[20]));
 sky130_fd_sc_hd__buf_12 output111 (.A(net111),
    .X(o_pc_IF[21]));
 sky130_fd_sc_hd__buf_12 output112 (.A(net112),
    .X(o_pc_IF[22]));
 sky130_fd_sc_hd__buf_12 output113 (.A(net113),
    .X(o_pc_IF[23]));
 sky130_fd_sc_hd__buf_12 output114 (.A(net114),
    .X(o_pc_IF[24]));
 sky130_fd_sc_hd__buf_12 output115 (.A(net115),
    .X(o_pc_IF[25]));
 sky130_fd_sc_hd__buf_12 output116 (.A(net116),
    .X(o_pc_IF[26]));
 sky130_fd_sc_hd__buf_12 output117 (.A(net117),
    .X(o_pc_IF[27]));
 sky130_fd_sc_hd__buf_12 output118 (.A(net118),
    .X(o_pc_IF[28]));
 sky130_fd_sc_hd__buf_12 output119 (.A(net119),
    .X(o_pc_IF[29]));
 sky130_fd_sc_hd__buf_12 output120 (.A(net120),
    .X(o_pc_IF[2]));
 sky130_fd_sc_hd__buf_12 output121 (.A(net121),
    .X(o_pc_IF[30]));
 sky130_fd_sc_hd__buf_12 output122 (.A(net122),
    .X(o_pc_IF[31]));
 sky130_fd_sc_hd__buf_12 output123 (.A(net123),
    .X(o_pc_IF[3]));
 sky130_fd_sc_hd__buf_12 output124 (.A(net124),
    .X(o_pc_IF[4]));
 sky130_fd_sc_hd__buf_12 output125 (.A(net125),
    .X(o_pc_IF[5]));
 sky130_fd_sc_hd__buf_12 output126 (.A(net126),
    .X(o_pc_IF[6]));
 sky130_fd_sc_hd__buf_12 output127 (.A(net127),
    .X(o_pc_IF[7]));
 sky130_fd_sc_hd__buf_12 output128 (.A(net128),
    .X(o_pc_IF[8]));
 sky130_fd_sc_hd__buf_12 output129 (.A(net129),
    .X(o_pc_IF[9]));
 sky130_fd_sc_hd__buf_12 output130 (.A(net130),
    .X(o_write_data_M[0]));
 sky130_fd_sc_hd__buf_12 output131 (.A(net131),
    .X(o_write_data_M[10]));
 sky130_fd_sc_hd__buf_12 output132 (.A(net132),
    .X(o_write_data_M[11]));
 sky130_fd_sc_hd__buf_12 output133 (.A(net133),
    .X(o_write_data_M[12]));
 sky130_fd_sc_hd__buf_12 output134 (.A(net134),
    .X(o_write_data_M[13]));
 sky130_fd_sc_hd__buf_12 output135 (.A(net135),
    .X(o_write_data_M[14]));
 sky130_fd_sc_hd__buf_12 output136 (.A(net136),
    .X(o_write_data_M[15]));
 sky130_fd_sc_hd__buf_12 output137 (.A(net137),
    .X(o_write_data_M[16]));
 sky130_fd_sc_hd__buf_12 output138 (.A(net138),
    .X(o_write_data_M[17]));
 sky130_fd_sc_hd__buf_12 output139 (.A(net139),
    .X(o_write_data_M[18]));
 sky130_fd_sc_hd__buf_12 output140 (.A(net140),
    .X(o_write_data_M[19]));
 sky130_fd_sc_hd__buf_12 output141 (.A(net141),
    .X(o_write_data_M[1]));
 sky130_fd_sc_hd__buf_12 output142 (.A(net142),
    .X(o_write_data_M[20]));
 sky130_fd_sc_hd__buf_12 output143 (.A(net143),
    .X(o_write_data_M[21]));
 sky130_fd_sc_hd__buf_12 output144 (.A(net144),
    .X(o_write_data_M[22]));
 sky130_fd_sc_hd__buf_12 output145 (.A(net145),
    .X(o_write_data_M[23]));
 sky130_fd_sc_hd__buf_12 output146 (.A(net146),
    .X(o_write_data_M[24]));
 sky130_fd_sc_hd__buf_12 output147 (.A(net147),
    .X(o_write_data_M[25]));
 sky130_fd_sc_hd__buf_12 output148 (.A(net148),
    .X(o_write_data_M[26]));
 sky130_fd_sc_hd__buf_12 output149 (.A(net149),
    .X(o_write_data_M[27]));
 sky130_fd_sc_hd__buf_12 output150 (.A(net150),
    .X(o_write_data_M[28]));
 sky130_fd_sc_hd__buf_12 output151 (.A(net151),
    .X(o_write_data_M[29]));
 sky130_fd_sc_hd__buf_12 output152 (.A(net152),
    .X(o_write_data_M[2]));
 sky130_fd_sc_hd__buf_12 output153 (.A(net153),
    .X(o_write_data_M[30]));
 sky130_fd_sc_hd__buf_12 output154 (.A(net154),
    .X(o_write_data_M[31]));
 sky130_fd_sc_hd__buf_12 output155 (.A(net155),
    .X(o_write_data_M[3]));
 sky130_fd_sc_hd__buf_12 output156 (.A(net156),
    .X(o_write_data_M[4]));
 sky130_fd_sc_hd__buf_12 output157 (.A(net157),
    .X(o_write_data_M[5]));
 sky130_fd_sc_hd__buf_12 output158 (.A(net158),
    .X(o_write_data_M[6]));
 sky130_fd_sc_hd__buf_12 output159 (.A(net159),
    .X(o_write_data_M[7]));
 sky130_fd_sc_hd__buf_12 output160 (.A(net160),
    .X(o_write_data_M[8]));
 sky130_fd_sc_hd__buf_12 output161 (.A(net161),
    .X(o_write_data_M[9]));
 sky130_fd_sc_hd__buf_12 output64 (.A(net64),
    .X(o_data_addr_M[0]));
 sky130_fd_sc_hd__buf_12 output65 (.A(net65),
    .X(o_data_addr_M[10]));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(o_data_addr_M[11]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(o_data_addr_M[12]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(o_data_addr_M[13]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(o_data_addr_M[14]));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(o_data_addr_M[15]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(o_data_addr_M[16]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net72),
    .X(o_data_addr_M[17]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(o_data_addr_M[18]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(o_data_addr_M[19]));
 sky130_fd_sc_hd__buf_12 output75 (.A(net75),
    .X(o_data_addr_M[1]));
 sky130_fd_sc_hd__buf_12 output76 (.A(net76),
    .X(o_data_addr_M[20]));
 sky130_fd_sc_hd__buf_12 output77 (.A(net77),
    .X(o_data_addr_M[21]));
 sky130_fd_sc_hd__buf_12 output78 (.A(net78),
    .X(o_data_addr_M[22]));
 sky130_fd_sc_hd__buf_12 output79 (.A(net79),
    .X(o_data_addr_M[23]));
 sky130_fd_sc_hd__buf_12 output80 (.A(net80),
    .X(o_data_addr_M[24]));
 sky130_fd_sc_hd__buf_12 output81 (.A(net81),
    .X(o_data_addr_M[25]));
 sky130_fd_sc_hd__buf_12 output82 (.A(net82),
    .X(o_data_addr_M[26]));
 sky130_fd_sc_hd__buf_12 output83 (.A(net83),
    .X(o_data_addr_M[27]));
 sky130_fd_sc_hd__buf_12 output84 (.A(net84),
    .X(o_data_addr_M[28]));
 sky130_fd_sc_hd__buf_12 output85 (.A(net85),
    .X(o_data_addr_M[29]));
 sky130_fd_sc_hd__buf_12 output86 (.A(net86),
    .X(o_data_addr_M[2]));
 sky130_fd_sc_hd__buf_12 output87 (.A(net87),
    .X(o_data_addr_M[30]));
 sky130_fd_sc_hd__buf_12 output88 (.A(net88),
    .X(o_data_addr_M[31]));
 sky130_fd_sc_hd__buf_12 output89 (.A(net89),
    .X(o_data_addr_M[3]));
 sky130_fd_sc_hd__buf_12 output90 (.A(net90),
    .X(o_data_addr_M[4]));
 sky130_fd_sc_hd__buf_12 output91 (.A(net91),
    .X(o_data_addr_M[5]));
 sky130_fd_sc_hd__buf_12 output92 (.A(net92),
    .X(o_data_addr_M[6]));
 sky130_fd_sc_hd__buf_12 output93 (.A(net93),
    .X(o_data_addr_M[7]));
 sky130_fd_sc_hd__buf_12 output94 (.A(net94),
    .X(o_data_addr_M[8]));
 sky130_fd_sc_hd__buf_12 output95 (.A(net95),
    .X(o_data_addr_M[9]));
 sky130_fd_sc_hd__buf_12 output96 (.A(net96),
    .X(o_funct3_MEM[0]));
 sky130_fd_sc_hd__buf_12 output97 (.A(net97),
    .X(o_funct3_MEM[1]));
 sky130_fd_sc_hd__buf_12 output98 (.A(net98),
    .X(o_funct3_MEM[2]));
 sky130_fd_sc_hd__buf_12 output99 (.A(net99),
    .X(o_mem_write_M));
 sky130_fd_sc_hd__buf_4 wire301 (.A(_2075_),
    .X(net301));
 assign o_pc_IF[0] = net476;
 assign o_pc_IF[1] = net477;
endmodule

