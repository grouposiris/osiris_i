// This is the unpowered netlist.
module osiris_i_mem (wb_clk_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input [4:0] io_in;
 output [6:0] io_oeb;
 output [1:0] io_out;

 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire \core_data_addr_M[0] ;
 wire \core_data_addr_M[10] ;
 wire \core_data_addr_M[11] ;
 wire \core_data_addr_M[12] ;
 wire \core_data_addr_M[13] ;
 wire \core_data_addr_M[14] ;
 wire \core_data_addr_M[15] ;
 wire \core_data_addr_M[16] ;
 wire \core_data_addr_M[17] ;
 wire \core_data_addr_M[18] ;
 wire \core_data_addr_M[19] ;
 wire \core_data_addr_M[1] ;
 wire \core_data_addr_M[20] ;
 wire \core_data_addr_M[21] ;
 wire \core_data_addr_M[22] ;
 wire \core_data_addr_M[23] ;
 wire \core_data_addr_M[24] ;
 wire \core_data_addr_M[25] ;
 wire \core_data_addr_M[26] ;
 wire \core_data_addr_M[27] ;
 wire \core_data_addr_M[28] ;
 wire \core_data_addr_M[29] ;
 wire \core_data_addr_M[2] ;
 wire \core_data_addr_M[30] ;
 wire \core_data_addr_M[31] ;
 wire \core_data_addr_M[3] ;
 wire \core_data_addr_M[4] ;
 wire \core_data_addr_M[5] ;
 wire \core_data_addr_M[6] ;
 wire \core_data_addr_M[7] ;
 wire \core_data_addr_M[8] ;
 wire \core_data_addr_M[9] ;
 wire \core_instr_ID[0] ;
 wire \core_instr_ID[10] ;
 wire \core_instr_ID[11] ;
 wire \core_instr_ID[12] ;
 wire \core_instr_ID[13] ;
 wire \core_instr_ID[14] ;
 wire \core_instr_ID[15] ;
 wire \core_instr_ID[16] ;
 wire \core_instr_ID[17] ;
 wire \core_instr_ID[18] ;
 wire \core_instr_ID[19] ;
 wire \core_instr_ID[1] ;
 wire \core_instr_ID[20] ;
 wire \core_instr_ID[21] ;
 wire \core_instr_ID[22] ;
 wire \core_instr_ID[23] ;
 wire \core_instr_ID[24] ;
 wire \core_instr_ID[25] ;
 wire \core_instr_ID[26] ;
 wire \core_instr_ID[27] ;
 wire \core_instr_ID[28] ;
 wire \core_instr_ID[29] ;
 wire \core_instr_ID[2] ;
 wire \core_instr_ID[30] ;
 wire \core_instr_ID[31] ;
 wire \core_instr_ID[3] ;
 wire \core_instr_ID[4] ;
 wire \core_instr_ID[5] ;
 wire \core_instr_ID[6] ;
 wire \core_instr_ID[7] ;
 wire \core_instr_ID[8] ;
 wire \core_instr_ID[9] ;
 wire core_mem_write_M;
 wire \core_pc_IF[0] ;
 wire \core_pc_IF[10] ;
 wire \core_pc_IF[11] ;
 wire \core_pc_IF[12] ;
 wire \core_pc_IF[13] ;
 wire \core_pc_IF[14] ;
 wire \core_pc_IF[15] ;
 wire \core_pc_IF[16] ;
 wire \core_pc_IF[17] ;
 wire \core_pc_IF[18] ;
 wire \core_pc_IF[19] ;
 wire \core_pc_IF[1] ;
 wire \core_pc_IF[20] ;
 wire \core_pc_IF[21] ;
 wire \core_pc_IF[22] ;
 wire \core_pc_IF[23] ;
 wire \core_pc_IF[24] ;
 wire \core_pc_IF[25] ;
 wire \core_pc_IF[26] ;
 wire \core_pc_IF[27] ;
 wire \core_pc_IF[28] ;
 wire \core_pc_IF[29] ;
 wire \core_pc_IF[2] ;
 wire \core_pc_IF[30] ;
 wire \core_pc_IF[31] ;
 wire \core_pc_IF[3] ;
 wire \core_pc_IF[4] ;
 wire \core_pc_IF[5] ;
 wire \core_pc_IF[6] ;
 wire \core_pc_IF[7] ;
 wire \core_pc_IF[8] ;
 wire \core_pc_IF[9] ;
 wire \core_read_data_M[0] ;
 wire \core_read_data_M[10] ;
 wire \core_read_data_M[11] ;
 wire \core_read_data_M[12] ;
 wire \core_read_data_M[13] ;
 wire \core_read_data_M[14] ;
 wire \core_read_data_M[15] ;
 wire \core_read_data_M[16] ;
 wire \core_read_data_M[17] ;
 wire \core_read_data_M[18] ;
 wire \core_read_data_M[19] ;
 wire \core_read_data_M[1] ;
 wire \core_read_data_M[20] ;
 wire \core_read_data_M[21] ;
 wire \core_read_data_M[22] ;
 wire \core_read_data_M[23] ;
 wire \core_read_data_M[24] ;
 wire \core_read_data_M[25] ;
 wire \core_read_data_M[26] ;
 wire \core_read_data_M[27] ;
 wire \core_read_data_M[28] ;
 wire \core_read_data_M[29] ;
 wire \core_read_data_M[2] ;
 wire \core_read_data_M[30] ;
 wire \core_read_data_M[31] ;
 wire \core_read_data_M[3] ;
 wire \core_read_data_M[4] ;
 wire \core_read_data_M[5] ;
 wire \core_read_data_M[6] ;
 wire \core_read_data_M[7] ;
 wire \core_read_data_M[8] ;
 wire \core_read_data_M[9] ;
 wire \core_write_data_M[0] ;
 wire \core_write_data_M[10] ;
 wire \core_write_data_M[11] ;
 wire \core_write_data_M[12] ;
 wire \core_write_data_M[13] ;
 wire \core_write_data_M[14] ;
 wire \core_write_data_M[15] ;
 wire \core_write_data_M[16] ;
 wire \core_write_data_M[17] ;
 wire \core_write_data_M[18] ;
 wire \core_write_data_M[19] ;
 wire \core_write_data_M[1] ;
 wire \core_write_data_M[20] ;
 wire \core_write_data_M[21] ;
 wire \core_write_data_M[22] ;
 wire \core_write_data_M[23] ;
 wire \core_write_data_M[24] ;
 wire \core_write_data_M[25] ;
 wire \core_write_data_M[26] ;
 wire \core_write_data_M[27] ;
 wire \core_write_data_M[28] ;
 wire \core_write_data_M[29] ;
 wire \core_write_data_M[2] ;
 wire \core_write_data_M[30] ;
 wire \core_write_data_M[31] ;
 wire \core_write_data_M[3] ;
 wire \core_write_data_M[4] ;
 wire \core_write_data_M[5] ;
 wire \core_write_data_M[6] ;
 wire \core_write_data_M[7] ;
 wire \core_write_data_M[8] ;
 wire \core_write_data_M[9] ;
 wire \data_mem_adr_i[2] ;
 wire \data_mem_adr_i[3] ;
 wire \data_mem_adr_i[4] ;
 wire \data_mem_adr_i[5] ;
 wire \data_mem_adr_i[6] ;
 wire \data_mem_adr_i[7] ;
 wire \data_reg[10] ;
 wire \data_reg[11] ;
 wire \data_reg[12] ;
 wire \data_reg[13] ;
 wire \data_reg[14] ;
 wire \data_reg[15] ;
 wire \data_reg[16] ;
 wire \data_reg[17] ;
 wire \data_reg[18] ;
 wire \data_reg[19] ;
 wire \data_reg[20] ;
 wire \data_reg[21] ;
 wire \data_reg[22] ;
 wire \data_reg[23] ;
 wire \data_reg[24] ;
 wire \data_reg[25] ;
 wire \data_reg[26] ;
 wire \data_reg[27] ;
 wire \data_reg[28] ;
 wire \data_reg[29] ;
 wire \data_reg[30] ;
 wire \data_reg[31] ;
 wire \data_reg[8] ;
 wire \data_reg[9] ;
 wire \dummy_data2[0] ;
 wire \dummy_data2[10] ;
 wire \dummy_data2[11] ;
 wire \dummy_data2[12] ;
 wire \dummy_data2[13] ;
 wire \dummy_data2[14] ;
 wire \dummy_data2[15] ;
 wire \dummy_data2[16] ;
 wire \dummy_data2[17] ;
 wire \dummy_data2[18] ;
 wire \dummy_data2[19] ;
 wire \dummy_data2[1] ;
 wire \dummy_data2[20] ;
 wire \dummy_data2[21] ;
 wire \dummy_data2[22] ;
 wire \dummy_data2[23] ;
 wire \dummy_data2[24] ;
 wire \dummy_data2[25] ;
 wire \dummy_data2[26] ;
 wire \dummy_data2[27] ;
 wire \dummy_data2[28] ;
 wire \dummy_data2[29] ;
 wire \dummy_data2[2] ;
 wire \dummy_data2[30] ;
 wire \dummy_data2[31] ;
 wire \dummy_data2[3] ;
 wire \dummy_data2[4] ;
 wire \dummy_data2[5] ;
 wire \dummy_data2[6] ;
 wire \dummy_data2[7] ;
 wire \dummy_data2[8] ;
 wire \dummy_data2[9] ;
 wire \dummy_data[0] ;
 wire \dummy_data[10] ;
 wire \dummy_data[11] ;
 wire \dummy_data[12] ;
 wire \dummy_data[13] ;
 wire \dummy_data[14] ;
 wire \dummy_data[15] ;
 wire \dummy_data[16] ;
 wire \dummy_data[17] ;
 wire \dummy_data[18] ;
 wire \dummy_data[19] ;
 wire \dummy_data[1] ;
 wire \dummy_data[20] ;
 wire \dummy_data[21] ;
 wire \dummy_data[22] ;
 wire \dummy_data[23] ;
 wire \dummy_data[24] ;
 wire \dummy_data[25] ;
 wire \dummy_data[26] ;
 wire \dummy_data[27] ;
 wire \dummy_data[28] ;
 wire \dummy_data[29] ;
 wire \dummy_data[2] ;
 wire \dummy_data[30] ;
 wire \dummy_data[31] ;
 wire \dummy_data[3] ;
 wire \dummy_data[4] ;
 wire \dummy_data[5] ;
 wire \dummy_data[6] ;
 wire \dummy_data[7] ;
 wire \dummy_data[8] ;
 wire \dummy_data[9] ;
 wire \funct3[0] ;
 wire \funct3[1] ;
 wire \funct3[2] ;
 wire \funct3_s2[0] ;
 wire \funct3_s2[1] ;
 wire \funct3_s2[2] ;
 wire \inst_mem_adr_i[0] ;
 wire \inst_mem_adr_i[1] ;
 wire \inst_mem_adr_i[2] ;
 wire \inst_mem_adr_i[3] ;
 wire \inst_mem_adr_i[4] ;
 wire \inst_mem_adr_i[5] ;
 wire \inst_mem_adr_i[6] ;
 wire \inst_mem_adr_i[7] ;
 wire \inst_mem_dat_i[0] ;
 wire \inst_mem_dat_i[10] ;
 wire \inst_mem_dat_i[11] ;
 wire \inst_mem_dat_i[12] ;
 wire \inst_mem_dat_i[13] ;
 wire \inst_mem_dat_i[14] ;
 wire \inst_mem_dat_i[15] ;
 wire \inst_mem_dat_i[16] ;
 wire \inst_mem_dat_i[17] ;
 wire \inst_mem_dat_i[18] ;
 wire \inst_mem_dat_i[19] ;
 wire \inst_mem_dat_i[1] ;
 wire \inst_mem_dat_i[20] ;
 wire \inst_mem_dat_i[21] ;
 wire \inst_mem_dat_i[22] ;
 wire \inst_mem_dat_i[23] ;
 wire \inst_mem_dat_i[24] ;
 wire \inst_mem_dat_i[25] ;
 wire \inst_mem_dat_i[26] ;
 wire \inst_mem_dat_i[27] ;
 wire \inst_mem_dat_i[28] ;
 wire \inst_mem_dat_i[29] ;
 wire \inst_mem_dat_i[2] ;
 wire \inst_mem_dat_i[30] ;
 wire \inst_mem_dat_i[31] ;
 wire \inst_mem_dat_i[3] ;
 wire \inst_mem_dat_i[4] ;
 wire \inst_mem_dat_i[5] ;
 wire \inst_mem_dat_i[6] ;
 wire \inst_mem_dat_i[7] ;
 wire \inst_mem_dat_i[8] ;
 wire \inst_mem_dat_i[9] ;
 wire \mux_funct3[0] ;
 wire \mux_funct3[1] ;
 wire \mux_funct3[2] ;
 wire \mux_funct3[3] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net32;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net394;
 wire net396;
 wire net397;
 wire net399;
 wire net4;
 wire net40;
 wire net401;
 wire net403;
 wire net41;
 wire net416;
 wire net418;
 wire net419;
 wire net42;
 wire net423;
 wire net43;
 wire net433;
 wire net438;
 wire net44;
 wire net441;
 wire net45;
 wire net451;
 wire net454;
 wire net46;
 wire net460;
 wire net463;
 wire net466;
 wire net47;
 wire net479;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire o_uart_tx;
 wire \shifted_data[0] ;
 wire \shifted_data[10] ;
 wire \shifted_data[11] ;
 wire \shifted_data[12] ;
 wire \shifted_data[13] ;
 wire \shifted_data[14] ;
 wire \shifted_data[15] ;
 wire \shifted_data[16] ;
 wire \shifted_data[17] ;
 wire \shifted_data[18] ;
 wire \shifted_data[19] ;
 wire \shifted_data[1] ;
 wire \shifted_data[20] ;
 wire \shifted_data[21] ;
 wire \shifted_data[22] ;
 wire \shifted_data[23] ;
 wire \shifted_data[24] ;
 wire \shifted_data[25] ;
 wire \shifted_data[26] ;
 wire \shifted_data[27] ;
 wire \shifted_data[28] ;
 wire \shifted_data[29] ;
 wire \shifted_data[2] ;
 wire \shifted_data[30] ;
 wire \shifted_data[31] ;
 wire \shifted_data[3] ;
 wire \shifted_data[4] ;
 wire \shifted_data[5] ;
 wire \shifted_data[6] ;
 wire \shifted_data[7] ;
 wire \shifted_data[8] ;
 wire \shifted_data[9] ;
 wire \uart_wb_adr_o[0] ;
 wire \uart_wb_adr_o[1] ;
 wire \uart_wb_adr_o[2] ;
 wire \uart_wb_adr_o[3] ;
 wire \uart_wb_adr_o[4] ;
 wire \uart_wb_adr_o[5] ;
 wire \uart_wb_adr_o[6] ;
 wire \uart_wb_adr_o[7] ;
 wire uart_wb_cyc_o;
 wire \uart_wb_dat_i[0] ;
 wire \uart_wb_dat_i[10] ;
 wire \uart_wb_dat_i[11] ;
 wire \uart_wb_dat_i[12] ;
 wire \uart_wb_dat_i[13] ;
 wire \uart_wb_dat_i[14] ;
 wire \uart_wb_dat_i[15] ;
 wire \uart_wb_dat_i[16] ;
 wire \uart_wb_dat_i[17] ;
 wire \uart_wb_dat_i[18] ;
 wire \uart_wb_dat_i[19] ;
 wire \uart_wb_dat_i[1] ;
 wire \uart_wb_dat_i[20] ;
 wire \uart_wb_dat_i[21] ;
 wire \uart_wb_dat_i[22] ;
 wire \uart_wb_dat_i[23] ;
 wire \uart_wb_dat_i[24] ;
 wire \uart_wb_dat_i[25] ;
 wire \uart_wb_dat_i[26] ;
 wire \uart_wb_dat_i[27] ;
 wire \uart_wb_dat_i[28] ;
 wire \uart_wb_dat_i[29] ;
 wire \uart_wb_dat_i[2] ;
 wire \uart_wb_dat_i[30] ;
 wire \uart_wb_dat_i[31] ;
 wire \uart_wb_dat_i[3] ;
 wire \uart_wb_dat_i[4] ;
 wire \uart_wb_dat_i[5] ;
 wire \uart_wb_dat_i[6] ;
 wire \uart_wb_dat_i[7] ;
 wire \uart_wb_dat_i[8] ;
 wire \uart_wb_dat_i[9] ;
 wire uart_wb_stb_o;
 wire uart_wb_we_o;
 wire write_sram_data_mem;
 wire write_sram_inst_mem;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\core_data_addr_M[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\core_data_addr_M[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\core_data_addr_M[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\core_data_addr_M[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\core_data_addr_M[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\core_data_addr_M[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(\core_pc_IF[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(\core_pc_IF[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\core_data_addr_M[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\core_data_addr_M[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\core_data_addr_M[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\core_data_addr_M[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\core_data_addr_M[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\core_data_addr_M[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\core_data_addr_M[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\core_data_addr_M[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(\core_read_data_M[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(\core_read_data_M[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(\core_read_data_M[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(\core_write_data_M[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(\core_write_data_M[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\core_data_addr_M[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(\core_write_data_M[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(\core_write_data_M[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(\core_write_data_M[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(\core_write_data_M[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(\core_write_data_M[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(\core_write_data_M[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(\core_write_data_M[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(\core_write_data_M[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(\core_write_data_M[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(\core_write_data_M[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\core_data_addr_M[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(\core_write_data_M[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(\core_write_data_M[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(\core_write_data_M[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(\core_write_data_M[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(\core_write_data_M[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(\core_write_data_M[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(\core_write_data_M[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(\core_write_data_M[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(\core_write_data_M[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(\core_write_data_M[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\core_data_addr_M[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(\data_reg[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(\data_reg[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(\data_reg[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(\data_reg[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(\data_reg[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(\data_reg[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(\data_reg[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(\data_reg[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_341 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_342 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_343 (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_344 (.DIODE(\data_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_345 (.DIODE(\data_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_346 (.DIODE(\data_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_347 (.DIODE(\data_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_348 (.DIODE(\data_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_349 (.DIODE(\data_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_350 (.DIODE(\data_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_351 (.DIODE(\data_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_352 (.DIODE(\data_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_353 (.DIODE(\data_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_354 (.DIODE(\data_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_355 (.DIODE(\data_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_356 (.DIODE(\inst_mem_dat_i[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_357 (.DIODE(\inst_mem_dat_i[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_358 (.DIODE(\inst_mem_dat_i[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_359 (.DIODE(\inst_mem_dat_i[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_360 (.DIODE(\inst_mem_dat_i[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_361 (.DIODE(\inst_mem_dat_i[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_362 (.DIODE(\inst_mem_dat_i[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_363 (.DIODE(\inst_mem_dat_i[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_364 (.DIODE(\inst_mem_dat_i[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_365 (.DIODE(\inst_mem_dat_i[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_366 (.DIODE(\inst_mem_dat_i[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_367 (.DIODE(\mux_funct3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_368 (.DIODE(\mux_funct3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_369 (.DIODE(\mux_funct3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_370 (.DIODE(\mux_funct3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_371 (.DIODE(\mux_funct3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_372 (.DIODE(\mux_funct3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_373 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_374 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_375 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_376 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_377 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_378 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_379 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_380 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_381 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_382 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_383 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_384 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_385 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_386 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_387 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_388 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_389 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_390 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_391 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_392 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_393 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_394 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_395 (.DIODE(\uart_wb_adr_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_396 (.DIODE(\uart_wb_adr_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_397 (.DIODE(\uart_wb_adr_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_398 (.DIODE(\uart_wb_adr_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_399 (.DIODE(\uart_wb_dat_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\core_data_addr_M[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_400 (.DIODE(\uart_wb_dat_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_401 (.DIODE(\uart_wb_dat_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_402 (.DIODE(\uart_wb_dat_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_403 (.DIODE(\uart_wb_dat_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_404 (.DIODE(\uart_wb_dat_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_405 (.DIODE(\uart_wb_dat_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_406 (.DIODE(\uart_wb_dat_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_407 (.DIODE(\uart_wb_dat_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_408 (.DIODE(\uart_wb_dat_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_409 (.DIODE(\uart_wb_dat_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_410 (.DIODE(\uart_wb_dat_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_411 (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_412 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_413 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_414 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_415 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_416 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_417 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_418 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_419 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_420 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_421 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_422 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_423 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_424 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_425 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_426 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_427 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_428 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_429 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_430 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_431 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_432 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_433 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_434 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_435 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_436 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_437 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_438 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_439 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_440 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_441 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_442 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_443 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_444 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_445 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_446 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_447 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_448 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_449 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_450 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_451 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_452 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_453 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_454 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_455 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_456 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_457 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_458 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_459 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_460 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_461 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_462 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_463 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_464 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_465 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_466 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_467 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_468 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_469 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_470 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_471 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_472 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_473 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_474 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_475 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_476 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_477 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_478 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_479 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_480 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_481 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_482 (.DIODE(\core_write_data_M[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_483 (.DIODE(\core_write_data_M[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_484 (.DIODE(\core_write_data_M[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_485 (.DIODE(\core_write_data_M[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_486 (.DIODE(\core_write_data_M[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_487 (.DIODE(\core_write_data_M[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_488 (.DIODE(\mux_funct3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_489 (.DIODE(\mux_funct3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_490 (.DIODE(\mux_funct3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_491 (.DIODE(\mux_funct3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_492 (.DIODE(\mux_funct3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_493 (.DIODE(\mux_funct3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_494 (.DIODE(\mux_funct3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_495 (.DIODE(\mux_funct3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_496 (.DIODE(\mux_funct3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_497 (.DIODE(\mux_funct3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_498 (.DIODE(\mux_funct3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_499 (.DIODE(\mux_funct3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\core_data_addr_M[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_500 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_501 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_502 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_503 (.DIODE(\mux_funct3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_504 (.DIODE(\mux_funct3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_505 (.DIODE(\mux_funct3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_506 (.DIODE(\mux_funct3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_507 (.DIODE(\mux_funct3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_508 (.DIODE(\mux_funct3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\core_data_addr_M[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\core_data_addr_M[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\core_data_addr_M[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\core_data_addr_M[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_U_CORE_clk (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[0]  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[10]  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[12]  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[13]  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[14]  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[15]  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[16]  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[17]  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[19]  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[20]  (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[21]  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[22]  (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[23]  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[24]  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[26]  (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[27]  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[28]  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[29]  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[2]  (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[30]  (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[3]  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[5]  (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[6]  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[7]  (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_instr_ID[9]  (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[0]  (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[10]  (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[11]  (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[12]  (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[14]  (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[15]  (.DIODE(\data_reg[15] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[17]  (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[18]  (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[19]  (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[1]  (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[20]  (.DIODE(\data_reg[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[22]  (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[23]  (.DIODE(\data_reg[23] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[24]  (.DIODE(\data_reg[24] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[25]  (.DIODE(\data_reg[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[26]  (.DIODE(\data_reg[26] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[27]  (.DIODE(\data_reg[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[28]  (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[29]  (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[2]  (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[30]  (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[31]  (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[3]  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[4]  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[5]  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[6]  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[7]  (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[8]  (.DIODE(\data_reg[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_CORE_i_read_data_M[9]  (.DIODE(\data_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_U_CORE_rst (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_U_DATA_MEM_clk0 (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[0]  (.DIODE(\shifted_data[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[10]  (.DIODE(\shifted_data[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[11]  (.DIODE(\shifted_data[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[12]  (.DIODE(\shifted_data[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[13]  (.DIODE(\shifted_data[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[14]  (.DIODE(\shifted_data[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[15]  (.DIODE(\shifted_data[15] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[16]  (.DIODE(\shifted_data[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[17]  (.DIODE(\shifted_data[17] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[18]  (.DIODE(\shifted_data[18] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[19]  (.DIODE(\shifted_data[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[1]  (.DIODE(\shifted_data[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[20]  (.DIODE(\shifted_data[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[21]  (.DIODE(\shifted_data[21] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[22]  (.DIODE(\shifted_data[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[23]  (.DIODE(\shifted_data[23] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[24]  (.DIODE(\shifted_data[24] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[25]  (.DIODE(\shifted_data[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[26]  (.DIODE(\shifted_data[26] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[27]  (.DIODE(\shifted_data[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[28]  (.DIODE(\shifted_data[28] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[29]  (.DIODE(\shifted_data[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[2]  (.DIODE(\shifted_data[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[30]  (.DIODE(\shifted_data[30] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[31]  (.DIODE(\shifted_data[31] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[3]  (.DIODE(\shifted_data[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[4]  (.DIODE(\shifted_data[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[5]  (.DIODE(\shifted_data[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[6]  (.DIODE(\shifted_data[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[7]  (.DIODE(\shifted_data[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[8]  (.DIODE(\shifted_data[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_DATA_MEM_din0[9]  (.DIODE(\shifted_data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_U_DATA_MEM_web0 (.DIODE(write_sram_data_mem));
 sky130_fd_sc_hd__diode_2 ANTENNA_U_INST_MEM_clk0 (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[0]  (.DIODE(\inst_mem_dat_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[10]  (.DIODE(\inst_mem_dat_i[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[11]  (.DIODE(\inst_mem_dat_i[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[12]  (.DIODE(\inst_mem_dat_i[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[13]  (.DIODE(\inst_mem_dat_i[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[14]  (.DIODE(\inst_mem_dat_i[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[15]  (.DIODE(\inst_mem_dat_i[15] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[16]  (.DIODE(\inst_mem_dat_i[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[17]  (.DIODE(\inst_mem_dat_i[17] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[18]  (.DIODE(\inst_mem_dat_i[18] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[19]  (.DIODE(\inst_mem_dat_i[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[1]  (.DIODE(\inst_mem_dat_i[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[20]  (.DIODE(\inst_mem_dat_i[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[21]  (.DIODE(\inst_mem_dat_i[21] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[22]  (.DIODE(\inst_mem_dat_i[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[23]  (.DIODE(\inst_mem_dat_i[23] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[24]  (.DIODE(\inst_mem_dat_i[24] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[25]  (.DIODE(\inst_mem_dat_i[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[26]  (.DIODE(\inst_mem_dat_i[26] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[27]  (.DIODE(\inst_mem_dat_i[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[28]  (.DIODE(\inst_mem_dat_i[28] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[29]  (.DIODE(\inst_mem_dat_i[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[2]  (.DIODE(\inst_mem_dat_i[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[30]  (.DIODE(\inst_mem_dat_i[30] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[31]  (.DIODE(\inst_mem_dat_i[31] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[3]  (.DIODE(\inst_mem_dat_i[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[4]  (.DIODE(\inst_mem_dat_i[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[5]  (.DIODE(\inst_mem_dat_i[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[6]  (.DIODE(\inst_mem_dat_i[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[7]  (.DIODE(\inst_mem_dat_i[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[8]  (.DIODE(\inst_mem_dat_i[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_INST_MEM_din0[9]  (.DIODE(\inst_mem_dat_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_U_INST_MEM_web0 (.DIODE(write_sram_inst_mem));
 sky130_fd_sc_hd__diode_2 ANTENNA_U_UART_WB_BRIDGE_clk (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_U_UART_WB_BRIDGE_i_start_rx (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_U_UART_WB_BRIDGE_i_uart_rx (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_U_UART_WB_BRIDGE_rst (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[0]  (.DIODE(\uart_wb_dat_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[10]  (.DIODE(\uart_wb_dat_i[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[11]  (.DIODE(\uart_wb_dat_i[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[12]  (.DIODE(\uart_wb_dat_i[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[13]  (.DIODE(\uart_wb_dat_i[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[14]  (.DIODE(\uart_wb_dat_i[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[16]  (.DIODE(\uart_wb_dat_i[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[17]  (.DIODE(\uart_wb_dat_i[17] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[18]  (.DIODE(\uart_wb_dat_i[18] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[19]  (.DIODE(\uart_wb_dat_i[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[1]  (.DIODE(\uart_wb_dat_i[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[20]  (.DIODE(\uart_wb_dat_i[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[21]  (.DIODE(\uart_wb_dat_i[21] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[23]  (.DIODE(\uart_wb_dat_i[23] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[24]  (.DIODE(\uart_wb_dat_i[24] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[25]  (.DIODE(\uart_wb_dat_i[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[26]  (.DIODE(\uart_wb_dat_i[26] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[27]  (.DIODE(\uart_wb_dat_i[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[28]  (.DIODE(\uart_wb_dat_i[28] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[29]  (.DIODE(\uart_wb_dat_i[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[2]  (.DIODE(\uart_wb_dat_i[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[30]  (.DIODE(\uart_wb_dat_i[30] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[31]  (.DIODE(\uart_wb_dat_i[31] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[3]  (.DIODE(\uart_wb_dat_i[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[4]  (.DIODE(\uart_wb_dat_i[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[5]  (.DIODE(\uart_wb_dat_i[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[6]  (.DIODE(\uart_wb_dat_i[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_U_UART_WB_BRIDGE_wb_dat_i[8]  (.DIODE(\uart_wb_dat_i[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__105__A (.DIODE(uart_wb_we_o));
 sky130_fd_sc_hd__diode_2 ANTENNA__106__B (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__107__B (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__108__A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__109__A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__109__C_N (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__110__B1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__111__A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__111__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__111__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__112__A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__112__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__113__A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__113__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__113__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__114__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__114__B2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__115__A_N (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__115__B (.DIODE(uart_wb_stb_o));
 sky130_fd_sc_hd__diode_2 ANTENNA__116__A1 (.DIODE(\core_pc_IF[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__116__S (.DIODE(_006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__117__A1 (.DIODE(\core_pc_IF[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__117__S (.DIODE(_006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__118__A1 (.DIODE(\core_pc_IF[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__118__S (.DIODE(_006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__119__A0 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__119__A1 (.DIODE(\core_pc_IF[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__119__S (.DIODE(_006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__A0 (.DIODE(\uart_wb_adr_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__A1 (.DIODE(\core_pc_IF[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__S (.DIODE(_006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__A0 (.DIODE(\uart_wb_adr_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__A1 (.DIODE(\core_pc_IF[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__S (.DIODE(_006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__A0 (.DIODE(\uart_wb_adr_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__A1 (.DIODE(\core_pc_IF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__S (.DIODE(_006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__A0 (.DIODE(\uart_wb_adr_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__A1 (.DIODE(\core_pc_IF[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__S (.DIODE(_006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__124__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__124__B (.DIODE(uart_wb_stb_o));
 sky130_fd_sc_hd__diode_2 ANTENNA__125__A1 (.DIODE(\core_data_addr_M[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__125__S (.DIODE(_007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__A0 (.DIODE(\uart_wb_adr_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__A1 (.DIODE(\core_data_addr_M[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__S (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__127__A0 (.DIODE(\uart_wb_adr_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__127__A1 (.DIODE(\core_data_addr_M[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__127__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__128__A0 (.DIODE(\uart_wb_adr_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__128__A1 (.DIODE(\core_data_addr_M[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__128__S (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__129__A0 (.DIODE(\uart_wb_adr_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__129__A1 (.DIODE(\core_data_addr_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__129__S (.DIODE(_007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__130__A0 (.DIODE(\uart_wb_adr_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__130__A1 (.DIODE(\core_data_addr_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__130__S (.DIODE(_007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__131__A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__131__B (.DIODE(uart_wb_stb_o));
 sky130_fd_sc_hd__diode_2 ANTENNA__132__A1 (.DIODE(\core_data_addr_M[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__132__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__133__A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__133__B (.DIODE(uart_wb_stb_o));
 sky130_fd_sc_hd__diode_2 ANTENNA__134__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__135__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__135__A2 (.DIODE(uart_wb_cyc_o));
 sky130_fd_sc_hd__diode_2 ANTENNA__135__B1 (.DIODE(\funct3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__135__B2 (.DIODE(\funct3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__135__C1 (.DIODE(\funct3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__136__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__136__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__136__B1 (.DIODE(_012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__137__A (.DIODE(\funct3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__137__B (.DIODE(\funct3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__137__C_N (.DIODE(\funct3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__A (.DIODE(\funct3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__B (.DIODE(\funct3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__C_N (.DIODE(\funct3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__139__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__139__B (.DIODE(_013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__139__C (.DIODE(_014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__A2 (.DIODE(_015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__B1 (.DIODE(_012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__141__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__141__A2 (.DIODE(_013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__141__B1 (.DIODE(_014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__A_N (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__143__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__143__A2 (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__143__B1 (.DIODE(_017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__143__C1 (.DIODE(_012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__A2 (.DIODE(_013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__145__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__145__A2 (.DIODE(uart_wb_cyc_o));
 sky130_fd_sc_hd__diode_2 ANTENNA__145__B1 (.DIODE(\funct3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__145__C1 (.DIODE(\funct3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__146__A0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__146__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__146__S (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__147__A0 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__147__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__147__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__148__A0 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__148__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__148__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__149__A0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__149__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__149__S (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__150__A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__150__A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__150__S (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__151__A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__151__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__151__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__152__A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__152__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__152__S (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__153__A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__153__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__153__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__154__A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__154__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__154__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__155__A0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__155__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__155__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__156__A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__156__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__156__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__157__A0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__157__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__157__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__A0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__159__A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__159__A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__159__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__160__A0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__160__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__160__S (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__161__A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__161__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__161__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__162__A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__162__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__162__S (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__163__A0 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__163__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__163__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__164__A0 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__164__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__164__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__165__A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__165__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__165__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__166__A0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__166__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__166__S (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__167__A0 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__167__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__167__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__168__A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__168__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__168__S (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__169__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__169__A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__169__S (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__170__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__170__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__170__S (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__171__A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__171__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__171__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__172__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__172__A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__172__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__173__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__173__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__173__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__174__A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__174__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__174__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__175__A0 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__175__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__175__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__176__A0 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__176__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__176__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__177__A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__177__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__177__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__178__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__178__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__178__B1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__179__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__179__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__179__B1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__180__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__180__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__180__B1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__B1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__182__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__182__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__182__B1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__183__A1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__183__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__183__B1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__B1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__185__A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__185__A3 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__185__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__186__A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__186__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__186__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__187__A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__187__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__188__A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__188__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__188__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__189__A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__189__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__189__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__190__A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__190__A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__190__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__191__A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__191__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__191__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__194__A1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__194__A2 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__194__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__195__A1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__195__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__196__A1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__196__A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__196__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__A1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__B1 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__198__B (.DIODE(_006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__199__A0 (.DIODE(uart_wb_we_o));
 sky130_fd_sc_hd__diode_2 ANTENNA__199__A1 (.DIODE(core_mem_write_M));
 sky130_fd_sc_hd__diode_2 ANTENNA__199__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__200__A (.DIODE(_019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__201__A0 (.DIODE(\inst_mem_dat_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__201__A1 (.DIODE(\core_write_data_M[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__201__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__202__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__202__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__202__C (.DIODE(_020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__203__A0 (.DIODE(\inst_mem_dat_i[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__203__A1 (.DIODE(\core_write_data_M[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__203__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__204__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__204__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__204__C (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__205__A0 (.DIODE(\inst_mem_dat_i[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__205__A1 (.DIODE(\core_write_data_M[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__205__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__206__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__206__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__206__C (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__207__A0 (.DIODE(\inst_mem_dat_i[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__207__A1 (.DIODE(\core_write_data_M[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__207__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__208__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__208__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__208__C (.DIODE(_023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__209__A0 (.DIODE(\inst_mem_dat_i[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__209__A1 (.DIODE(\core_write_data_M[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__209__S (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__210__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__210__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__210__C (.DIODE(_024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__211__A0 (.DIODE(\inst_mem_dat_i[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__211__A1 (.DIODE(\core_write_data_M[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__211__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__212__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__212__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__212__C (.DIODE(_025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__213__A0 (.DIODE(\inst_mem_dat_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__213__A1 (.DIODE(\core_write_data_M[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__213__S (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__214__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__214__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__214__C (.DIODE(_026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__215__A0 (.DIODE(\inst_mem_dat_i[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__215__A1 (.DIODE(\core_write_data_M[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__215__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__216__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__216__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__216__C (.DIODE(_027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__217__A0 (.DIODE(\inst_mem_dat_i[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__217__A1 (.DIODE(\core_write_data_M[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__217__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__218__A0 (.DIODE(_020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__218__A1 (.DIODE(_028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__218__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__219__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__219__B (.DIODE(_029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__220__A0 (.DIODE(\inst_mem_dat_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__220__A1 (.DIODE(\core_write_data_M[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__220__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__221__A0 (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__221__A1 (.DIODE(_030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__221__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__222__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__222__B (.DIODE(_031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__223__A0 (.DIODE(\inst_mem_dat_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__223__A1 (.DIODE(\core_write_data_M[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__223__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__224__A0 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__224__A1 (.DIODE(_032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__224__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__225__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__225__B (.DIODE(_033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__226__A0 (.DIODE(\inst_mem_dat_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__226__A1 (.DIODE(\core_write_data_M[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__226__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__227__A0 (.DIODE(_023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__227__A1 (.DIODE(_034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__227__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__228__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__228__B (.DIODE(_035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__229__A0 (.DIODE(\inst_mem_dat_i[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__229__A1 (.DIODE(\core_write_data_M[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__229__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__230__A0 (.DIODE(_024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__230__A1 (.DIODE(_036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__230__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__231__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__231__B (.DIODE(_037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__232__A0 (.DIODE(\inst_mem_dat_i[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__232__A1 (.DIODE(\core_write_data_M[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__232__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__233__A0 (.DIODE(_025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__233__A1 (.DIODE(_038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__233__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__234__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__234__B (.DIODE(_039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__235__A0 (.DIODE(\inst_mem_dat_i[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__235__A1 (.DIODE(\core_write_data_M[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__235__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__236__A0 (.DIODE(_026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__236__A1 (.DIODE(_040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__236__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__237__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__237__B (.DIODE(_041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__238__A0 (.DIODE(\inst_mem_dat_i[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__238__A1 (.DIODE(\core_write_data_M[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__238__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__A0 (.DIODE(_027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__A1 (.DIODE(_042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__240__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__240__B (.DIODE(_043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__241__A0 (.DIODE(\inst_mem_dat_i[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__241__A1 (.DIODE(\core_write_data_M[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__241__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__242__A0 (.DIODE(_028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__242__A1 (.DIODE(_044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__242__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__A1 (.DIODE(_017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__A2 (.DIODE(_020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__B1 (.DIODE(_045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__244__A0 (.DIODE(\inst_mem_dat_i[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__244__A1 (.DIODE(\core_write_data_M[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__244__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__245__A0 (.DIODE(_030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__245__A1 (.DIODE(_046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__245__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__246__A1 (.DIODE(_017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__246__A2 (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__246__B1 (.DIODE(_047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__246__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__247__A0 (.DIODE(\inst_mem_dat_i[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__247__A1 (.DIODE(\core_write_data_M[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__247__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__248__A0 (.DIODE(_032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__248__A1 (.DIODE(_048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__248__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__249__A1 (.DIODE(_017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__249__A2 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__249__B1 (.DIODE(_049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__249__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__250__A0 (.DIODE(\inst_mem_dat_i[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__250__A1 (.DIODE(\core_write_data_M[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__250__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__251__A0 (.DIODE(_034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__251__A1 (.DIODE(_050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__251__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__252__A1 (.DIODE(_017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__252__A2 (.DIODE(_023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__252__B1 (.DIODE(_051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__252__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__253__A0 (.DIODE(\inst_mem_dat_i[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__253__A1 (.DIODE(\core_write_data_M[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__253__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__254__A0 (.DIODE(_036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__254__A1 (.DIODE(_052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__254__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__255__A1 (.DIODE(_017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__255__A2 (.DIODE(_024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__255__B1 (.DIODE(_053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__255__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__256__A0 (.DIODE(\inst_mem_dat_i[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__256__A1 (.DIODE(\core_write_data_M[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__256__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__257__A0 (.DIODE(_038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__257__A1 (.DIODE(_054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__257__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__A1 (.DIODE(_017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__A2 (.DIODE(_025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__B1 (.DIODE(_055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__B2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__259__A0 (.DIODE(\inst_mem_dat_i[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__259__A1 (.DIODE(\core_write_data_M[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__259__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__260__A0 (.DIODE(_040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__260__A1 (.DIODE(_056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__260__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__261__A1 (.DIODE(_017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__261__A2 (.DIODE(_026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__261__B1 (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__261__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__262__A0 (.DIODE(\inst_mem_dat_i[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__262__A1 (.DIODE(\core_write_data_M[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__262__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__263__A0 (.DIODE(_042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__263__A1 (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__263__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__A1 (.DIODE(_017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__A2 (.DIODE(_027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__B1 (.DIODE(_059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__B2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__265__A0 (.DIODE(\inst_mem_dat_i[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__265__A1 (.DIODE(\core_write_data_M[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__265__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__266__A0 (.DIODE(_044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__266__A1 (.DIODE(_060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__266__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__267__A0 (.DIODE(_029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__267__A1 (.DIODE(_061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__267__S (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__268__A0 (.DIODE(\inst_mem_dat_i[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__268__A1 (.DIODE(\core_write_data_M[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__268__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__269__A0 (.DIODE(_046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__269__A1 (.DIODE(_062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__269__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__270__A0 (.DIODE(_031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__270__A1 (.DIODE(_063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__270__S (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__271__A0 (.DIODE(\inst_mem_dat_i[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__271__A1 (.DIODE(\core_write_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__271__S (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__272__A0 (.DIODE(_048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__272__A1 (.DIODE(_064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__272__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__273__A0 (.DIODE(_033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__273__A1 (.DIODE(_065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__273__S (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__274__A0 (.DIODE(\inst_mem_dat_i[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__274__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__275__A0 (.DIODE(_050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__275__A1 (.DIODE(_066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__275__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__276__A0 (.DIODE(_035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__276__A1 (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__276__S (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__277__A0 (.DIODE(\inst_mem_dat_i[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__277__A1 (.DIODE(\core_write_data_M[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__277__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__278__A0 (.DIODE(_052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__278__A1 (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__278__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__279__A0 (.DIODE(_037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__279__A1 (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__279__S (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__280__A0 (.DIODE(\inst_mem_dat_i[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__280__A1 (.DIODE(\core_write_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__280__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__281__A0 (.DIODE(_054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__281__A1 (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__281__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__282__A0 (.DIODE(_039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__282__A1 (.DIODE(_071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__282__S (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__283__A0 (.DIODE(\inst_mem_dat_i[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__283__S (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__284__A0 (.DIODE(_056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__284__A1 (.DIODE(_072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__284__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__285__A0 (.DIODE(_041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__285__A1 (.DIODE(_073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__285__S (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__286__A0 (.DIODE(\inst_mem_dat_i[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__286__A1 (.DIODE(\core_write_data_M[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__286__S (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__287__A0 (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__287__A1 (.DIODE(_074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__287__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__288__A0 (.DIODE(_043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__288__A1 (.DIODE(_075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__288__S (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__289__CLK (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__289__D (.DIODE(\funct3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__290__CLK (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__290__D (.DIODE(\funct3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__291__CLK (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__291__D (.DIODE(\funct3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__328__A (.DIODE(o_uart_tx));
 sky130_fd_sc_hd__diode_2 ANTENNA__329__A (.DIODE(o_uart_tx));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout12_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout13_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout14_A (.DIODE(_011_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout15_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout16_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout17_A (.DIODE(_009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout19_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout20_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout21_A (.DIODE(_007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout22_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout311_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold103_A (.DIODE(\data_reg[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold117_A (.DIODE(\data_reg[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold120_A (.DIODE(\data_reg[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold132_A (.DIODE(\data_reg[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold51_A (.DIODE(\data_reg[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold5_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold63_A (.DIODE(\data_reg[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold72_A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold82_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold84_A (.DIODE(\data_reg[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold94_A (.DIODE(\data_reg[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold9_A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap115_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap121_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap127_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap151_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap177_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap18_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap27_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap280_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap285_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap289_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap33_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap40_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap47_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap53_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap58_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap68_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap78_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap83_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap99_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire101_A (.DIODE(\core_instr_ID[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire102_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire103_A (.DIODE(\core_instr_ID[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire104_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire105_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire108_A (.DIODE(\core_instr_ID[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire109_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire10_A (.DIODE(\mux_funct3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire110_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire112_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire113_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire114_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire116_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire117_A (.DIODE(\core_instr_ID[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire118_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire119_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire11_A (.DIODE(\mux_funct3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire120_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire122_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire124_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire125_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire126_A (.DIODE(\core_instr_ID[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire128_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire129_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire131_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire132_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire134_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire135_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire136_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire138_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire139_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire140_A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire142_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire144_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire145_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire147_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire148_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire149_A (.DIODE(\core_instr_ID[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire150_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire153_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire154_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire155_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire156_A (.DIODE(\core_read_data_M[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire157_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire158_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire159_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire161_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire162_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire163_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire164_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire166_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire167_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire168_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire171_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire173_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire174_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire176_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire178_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire179_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire180_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire182_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire183_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire184_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire185_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire187_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire190_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire191_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire193_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire196_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire197_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire199_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire200_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire201_A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire202_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire204_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire205_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire206_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire207_A (.DIODE(\core_read_data_M[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire208_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire211_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire212_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire214_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire216_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire217_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire219_A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire220_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire221_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire222_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire223_A (.DIODE(\core_read_data_M[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire225_A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire228_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire229_A (.DIODE(\core_read_data_M[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire230_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire232_A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire233_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire235_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire238_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire239_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire23_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire241_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire244_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire245_A (.DIODE(\core_read_data_M[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire246_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire248_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire249_A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire24_A (.DIODE(\core_instr_ID[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire251_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire253_A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire254_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire256_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire257_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire258_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire259_A (.DIODE(\core_read_data_M[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire25_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire260_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire263_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire265_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire267_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire268_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire270_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire272_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire273_A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire275_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire277_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire278_A (.DIODE(\core_read_data_M[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire282_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire286_A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire287_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire28_A (.DIODE(\core_instr_ID[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire290_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire291_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire293_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire294_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire295_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire297_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire298_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire299_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire29_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire301_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire302_A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire303_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire305_A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire306_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire307_A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire30_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire31_A (.DIODE(\core_instr_ID[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire32_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire34_A (.DIODE(\core_instr_ID[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire35_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire36_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire37_A (.DIODE(\core_instr_ID[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire38_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire41_A (.DIODE(\core_instr_ID[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire42_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire43_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire44_A (.DIODE(\core_instr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire45_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire48_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire49_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire50_A (.DIODE(\core_instr_ID[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire51_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire52_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire54_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire55_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire57_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire59_A (.DIODE(\core_instr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire60_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire61_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire62_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire63_A (.DIODE(\core_instr_ID[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire65_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire66_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire67_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire69_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire70_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire72_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire73_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire74_A (.DIODE(\core_instr_ID[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire75_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire76_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire77_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire79_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire80_A (.DIODE(\core_instr_ID[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire81_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire84_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire85_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire87_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire88_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire8_A (.DIODE(\mux_funct3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire90_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire91_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire92_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire93_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire95_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire96_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire98_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire9_A (.DIODE(\mux_funct3[2] ));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_2385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2010 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_2022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_2030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_2036 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_2038 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_2063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2078 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2094 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_2106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_2190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_2234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_2259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1822 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1924 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1926 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_2024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_2254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_2310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_2478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_2534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_2590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_2646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1942 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1954 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_2002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_2006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_2010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_2014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_2018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_2022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_2026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_2054 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_2282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_2338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_2562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_2568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1924 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_2018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_2024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_2254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_2310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_2478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_2534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_2590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_2646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_2058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_2246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_2254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_2259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_2263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_2267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_2274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_2278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_2286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_2562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_2031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_2242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_2282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_2306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_2478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_2534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_2590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_2646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1898 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_2243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_2286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_2614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_2026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_2186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_2196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_2206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_2229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_2310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_2363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_2480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_2484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_2554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_2557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_2565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_2570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_2576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_2587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_2594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_2602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_2606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1882 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1924 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1952 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_2006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_2010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_2025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2036 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_2059 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2078 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_2162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_2170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_2206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_2248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_2414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_2424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_2442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_2452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_2458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_2503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_2538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_2542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_2602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_2630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_2645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_2654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_2665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_2742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_2754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_2766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_2778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_2738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_2742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_2774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_2774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_2738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_2774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1784 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1730 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_2738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_2742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_2738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_2742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_2746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_2754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_2766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_2778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_2738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_2742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_2746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_2750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_2754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_2758 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_2760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_2766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_2743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_2747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_2751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_2755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_2759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_2763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_2767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_2775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_2738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_2742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_2746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_2750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_2754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_2760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_2764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_2768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_2738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_2742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_2750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_2768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_2780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_2738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1730 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1702 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_2760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_2772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_1809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_1774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_2774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_1745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_1717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_1801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_1762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_1785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_1677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_1721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_1725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_1661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_1706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_1803 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_1412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_1613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_1773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_1809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_2738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_1717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_1721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_1725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_2742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_2754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_2766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_2778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_1295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_1709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_1793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_2738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_2742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_2746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_2750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_2754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_2758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_2760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_2764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_2768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_2772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_1747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_1755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_1794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_1802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_2742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_2754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_2766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_2778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_1798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_1804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_1809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_1799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_2774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_2788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_2800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_1786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_1798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_1719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_1727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_1811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_1792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_1796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_1800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1756 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_1778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_1798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_1766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_1771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_1775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_1779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_1783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_1792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_1796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_1801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_1812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_2738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_1702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_1710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_1782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_1792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_2742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_2754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_2766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_2778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_1730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_1769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_1783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_1802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_2738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_2742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_2746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_2738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_2742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_2746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_2750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_2754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_2758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_2766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_2778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_1657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_1661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_1665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230_1669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230_1730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_1742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_1746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_1774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_2738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_2742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_1794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_231_1802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_2774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_232_1657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_1718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_232_1766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_1782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_232_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_232_1797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_1794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_233_1802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_2758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_2770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_2778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_2781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_1812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_2738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_2742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_2758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_2760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234_2768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_2773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_2777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_2781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_2789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_2801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_1747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_1755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_1794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_235_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_2740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_2751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_2755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_2759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_2763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_2767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_2771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_2775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_2781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_2785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_2788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_2792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_2796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_1794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_1798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_2738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_2760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_236_2772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_2777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_2781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_2789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_2801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_1796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_2758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_2770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_2778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_2781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238_1801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_2742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_238_2754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_1782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_1794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_1802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_242_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_1664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_242_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_1809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_244_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_1652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1784 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244_1795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_1803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_2742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_244_2754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_1648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_245_1654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_1669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_1673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_245_1782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_1802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_245_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_245_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_246_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_2742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_246_2754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_247_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_247_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_1686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_1708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_248_1809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_1787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_1791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_1795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_1809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_250_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1784 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250_1795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_250_1799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_251_1684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_251_1806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_251_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_251_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_251_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_251_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_252_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_252_1674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_252_1685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_252_1700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_252_1704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_252_1720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_252_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_252_1794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_252_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_254_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_254_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_255_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_255_1782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_255_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_255_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_255_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_255_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_256_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_256_1669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_256_1754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_256_1781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_256_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_256_1792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_256_1806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_256_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_256_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_2738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_256_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_257_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_257_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_257_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_258_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1784 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_258_1795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_258_1803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_259_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_259_1782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_259_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_259_1807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_259_1811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_259_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_259_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_259_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_260_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_260_1669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_260_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_260_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_261_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_261_1702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_261_1723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_261_1731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_261_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_261_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_261_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_261_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_262_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_262_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_262_1794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_262_1812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_263_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_263_1781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_263_1787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_263_1791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_263_1796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_263_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_263_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_263_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_263_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_264_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_264_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_264_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_265_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_265_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_265_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_265_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_265_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_265_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_266_1669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_266_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_266_1794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_266_1804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_266_1812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267_1656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_267_1794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_267_1799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267_1804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267_1808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_267_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_267_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_268_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_268_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268_1797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268_1808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268_1812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_269_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_269_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_269_1801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_269_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_269_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_269_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_269_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_270_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_270_1669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_270_1798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_271_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_271_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_271_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_271_1809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_271_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_271_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_271_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_272_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_272_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_272_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_272_1812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_273_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_273_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_273_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_273_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_273_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_273_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_274_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_274_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_274_1804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_274_1808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_275_1672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_1699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_275_1770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_1781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_1785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_1789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_1804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_1808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_275_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_275_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_276_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_276_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_276_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_277_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_277_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_277_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_277_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_277_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_278_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_279_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_279_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_279_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_279_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_279_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_280_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_280_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_280_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_280_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_2738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_280_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_281_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_282_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_282_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_283_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_283_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_283_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_283_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_284_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_284_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_285_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_285_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_285_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_285_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_285_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_286_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_286_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_286_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_286_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_287_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_287_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_287_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_287_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_288_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_288_1652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_288_1658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_288_1662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_288_1670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_288_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_289_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_289_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_289_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_2742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_2754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_2766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_289_2778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_289_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_289_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_290_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_290_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_290_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_291_1652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_291_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_291_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_291_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_291_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_291_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_292_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_292_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_292_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_292_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_293_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_293_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_293_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_293_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_294_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_294_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_294_1664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_294_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_295_1652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_295_1658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_295_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_295_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_295_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_295_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_296_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_296_1651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_296_1658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_296_1662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_296_1670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_296_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_297_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_297_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_297_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_297_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_297_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_298_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_298_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_298_1664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_298_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_299_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_300_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_300_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_301_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_301_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_301_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_301_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_302_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_302_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_303_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_303_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_303_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_303_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_304_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_304_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_304_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_2738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_304_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_305_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_305_1692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_305_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_305_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_305_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_306_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_306_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_306_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_307_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_307_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_307_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_307_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_308_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_308_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_308_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_308_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_310_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_310_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_311_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_311_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_311_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_311_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_312_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_312_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_313_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_313_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_313_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_313_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_313_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_314_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_314_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_314_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_2738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_314_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_315_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_315_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_315_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_315_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_316_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_316_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_316_1664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_316_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_317_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_317_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_317_1794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_317_1802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_317_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_317_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_317_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_318_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_318_1798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_319_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_319_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_319_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_319_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_319_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_320_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_320_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_320_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_320_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_322_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_322_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_323_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_323_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_323_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_323_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_324_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_324_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_1656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_324_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_324_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_325_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_325_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_325_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_325_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_326_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_326_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_327_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_2767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_327_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_327_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_327_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_328_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_328_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_329_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_329_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_329_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_329_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_330_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_330_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_331_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_332_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_332_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_333_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_333_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_333_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_333_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_334_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_334_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_335_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_335_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_335_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_335_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_336_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_336_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_337_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_337_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_337_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_338_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_338_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_338_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_2738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_338_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_339_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_339_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_339_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_339_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_340_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_340_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_341_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_341_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_341_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_341_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_342_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_342_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_343_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_343_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_343_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_343_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_344_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_344_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_2796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_344_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_345_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_345_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_345_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_345_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_346_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_1786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_346_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_346_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_346_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_2738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_346_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_347_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_347_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_347_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_347_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_348_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_348_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_1794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_349_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_2084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_2092 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_2094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_2100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_2103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_2119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_2122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_2128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_2131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_2139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_2148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_2168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_2252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_2260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_2262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_2287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_2302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_2310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_2313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_350_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_1786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_350_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_350_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_350_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_351_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_1782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_351_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_351_1801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_351_1805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_351_1809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_351_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_2774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_351_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_351_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_1786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_352_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_352_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_352_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_352_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_353_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_1794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_353_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_353_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_353_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_353_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_354_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_1786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_354_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_354_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_355_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_1782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_355_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_355_1801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_355_1805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_355_1809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_355_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_355_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_355_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_356_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_356_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_1652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_356_1664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_1786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_356_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_356_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_357_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_1794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_357_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_357_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_357_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_357_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_358_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_359_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_359_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_1664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_1688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_359_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_359_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_359_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_359_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_359_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_360_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_1651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_360_1663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_360_1671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_360_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_360_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_360_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_360_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_360_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_360_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_360_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_360_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_2742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_360_2754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_360_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_360_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_360_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_360_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_361_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_361_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_361_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_361_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_361_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_361_2738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_361_2742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_361_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_361_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_361_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_362_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_362_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_362_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_362_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_362_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_362_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_362_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_362_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_2742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_362_2754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_362_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_362_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_362_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_362_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_363_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_363_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_363_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_363_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_363_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_363_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_363_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_364_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_364_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_364_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_364_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_364_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_364_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_364_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_364_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_364_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_364_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_364_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_364_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_1794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_366_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_366_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_366_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_366_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_366_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_366_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_366_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_366_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_366_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_2738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_366_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_366_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_366_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_366_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_366_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_367_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_367_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_367_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_367_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_367_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_367_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_367_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_368_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_368_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_368_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_368_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_368_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_368_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_368_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_368_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_368_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_368_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_368_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_368_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_369_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_369_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_369_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_369_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_369_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_369_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_2742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_2754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_2766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_369_2778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_369_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_369_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_370_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_370_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_370_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_370_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_370_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_370_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_370_1810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_370_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_370_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_370_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_370_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_370_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_370_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_371_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_371_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_371_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_371_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_371_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_371_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_371_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_372_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_1648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_372_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_372_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_372_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_372_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_372_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_372_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_372_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_372_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_372_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_372_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_372_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_372_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_373_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_373_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_373_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_373_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_2746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_373_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373_2786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_2788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_2800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_373_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_373_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_374_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_374_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_374_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_374_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_374_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_374_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_1798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_374_1810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_374_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_2746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_374_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_2772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_2784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_374_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_374_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_374_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_1838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375_1858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375_1864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_1966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_1978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375_1982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_1986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_1989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_1993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_1997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375_2010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_2014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375_2033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2038 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375_2042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_2046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_375_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_375_2078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_2086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_375_2110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375_2134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375_2200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_2204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_375_2222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_375_2250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_375_2306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_375_2318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_2344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_375_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_375_2414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375_2424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375_2514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_2518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_375_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375_2570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_2574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_375_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_375_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_2658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_375_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_375_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_375_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_376_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_1946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_1966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_376_1978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_1986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_376_1989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_376_1993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_376_1997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_376_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_376_2049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_2090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_376_2098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_2282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_376_2326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_376_2336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_376_2514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_376_2525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_376_2565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_376_2570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_376_2577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_376_2581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_376_2585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_376_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_377_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_1974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_1980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_377_1982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_1990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_1993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_377_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_2086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_2142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_2254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_2260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_2310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_2316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_2422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_2478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_2534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_2540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_2590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_2596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_2646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_2702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_2758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_2764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_2802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_377_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_378_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_1946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_1990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_378_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_379_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_379_1299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_379_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_1355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_1367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_379_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_1422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_379_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_379_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_379_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_379_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_379_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_379_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_379_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_380_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_380_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_380_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_380_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_380_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_380_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_380_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_380_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_380_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_380_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_380_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_380_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_380_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_380_1380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_380_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_380_1391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_380_1402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_380_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_380_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_380_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_380_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_380_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_380_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_380_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_380_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_381_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_381_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_381_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_381_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_381_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_381_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_381_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_381_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_381_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_381_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_382_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_383_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_384_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_385_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_386_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_387_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_388_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_389_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_390_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_391_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_392_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_394_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_395_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_396_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_397_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_398_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_399_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_2369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_2373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_2413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_400_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_401_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_401_1839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_401_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_401_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_401_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_401_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_2369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_2373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_2377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_2381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_2385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1924 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_2369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_2373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_2413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1924 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1926 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_2385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1924 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_2385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1924 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1924 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_2443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_2779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_2811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_2795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_2807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_989 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_1000 ();
 sky130_fd_sc_hd__decap_3 PHY_1001 ();
 sky130_fd_sc_hd__decap_3 PHY_1002 ();
 sky130_fd_sc_hd__decap_3 PHY_1003 ();
 sky130_fd_sc_hd__decap_3 PHY_1004 ();
 sky130_fd_sc_hd__decap_3 PHY_1005 ();
 sky130_fd_sc_hd__decap_3 PHY_1006 ();
 sky130_fd_sc_hd__decap_3 PHY_1007 ();
 sky130_fd_sc_hd__decap_3 PHY_1008 ();
 sky130_fd_sc_hd__decap_3 PHY_1009 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_1010 ();
 sky130_fd_sc_hd__decap_3 PHY_1011 ();
 sky130_fd_sc_hd__decap_3 PHY_1012 ();
 sky130_fd_sc_hd__decap_3 PHY_1013 ();
 sky130_fd_sc_hd__decap_3 PHY_1014 ();
 sky130_fd_sc_hd__decap_3 PHY_1015 ();
 sky130_fd_sc_hd__decap_3 PHY_1016 ();
 sky130_fd_sc_hd__decap_3 PHY_1017 ();
 sky130_fd_sc_hd__decap_3 PHY_1018 ();
 sky130_fd_sc_hd__decap_3 PHY_1019 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_1020 ();
 sky130_fd_sc_hd__decap_3 PHY_1021 ();
 sky130_fd_sc_hd__decap_3 PHY_1022 ();
 sky130_fd_sc_hd__decap_3 PHY_1023 ();
 sky130_fd_sc_hd__decap_3 PHY_1024 ();
 sky130_fd_sc_hd__decap_3 PHY_1025 ();
 sky130_fd_sc_hd__decap_3 PHY_1026 ();
 sky130_fd_sc_hd__decap_3 PHY_1027 ();
 sky130_fd_sc_hd__decap_3 PHY_1028 ();
 sky130_fd_sc_hd__decap_3 PHY_1029 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_1030 ();
 sky130_fd_sc_hd__decap_3 PHY_1031 ();
 sky130_fd_sc_hd__decap_3 PHY_1032 ();
 sky130_fd_sc_hd__decap_3 PHY_1033 ();
 sky130_fd_sc_hd__decap_3 PHY_1034 ();
 sky130_fd_sc_hd__decap_3 PHY_1035 ();
 sky130_fd_sc_hd__decap_3 PHY_1036 ();
 sky130_fd_sc_hd__decap_3 PHY_1037 ();
 sky130_fd_sc_hd__decap_3 PHY_1038 ();
 sky130_fd_sc_hd__decap_3 PHY_1039 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_1040 ();
 sky130_fd_sc_hd__decap_3 PHY_1041 ();
 sky130_fd_sc_hd__decap_3 PHY_1042 ();
 sky130_fd_sc_hd__decap_3 PHY_1043 ();
 sky130_fd_sc_hd__decap_3 PHY_1044 ();
 sky130_fd_sc_hd__decap_3 PHY_1045 ();
 sky130_fd_sc_hd__decap_3 PHY_1046 ();
 sky130_fd_sc_hd__decap_3 PHY_1047 ();
 sky130_fd_sc_hd__decap_3 PHY_1048 ();
 sky130_fd_sc_hd__decap_3 PHY_1049 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_1050 ();
 sky130_fd_sc_hd__decap_3 PHY_1051 ();
 sky130_fd_sc_hd__decap_3 PHY_1052 ();
 sky130_fd_sc_hd__decap_3 PHY_1053 ();
 sky130_fd_sc_hd__decap_3 PHY_1054 ();
 sky130_fd_sc_hd__decap_3 PHY_1055 ();
 sky130_fd_sc_hd__decap_3 PHY_1056 ();
 sky130_fd_sc_hd__decap_3 PHY_1057 ();
 sky130_fd_sc_hd__decap_3 PHY_1058 ();
 sky130_fd_sc_hd__decap_3 PHY_1059 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_1060 ();
 sky130_fd_sc_hd__decap_3 PHY_1061 ();
 sky130_fd_sc_hd__decap_3 PHY_1062 ();
 sky130_fd_sc_hd__decap_3 PHY_1063 ();
 sky130_fd_sc_hd__decap_3 PHY_1064 ();
 sky130_fd_sc_hd__decap_3 PHY_1065 ();
 sky130_fd_sc_hd__decap_3 PHY_1066 ();
 sky130_fd_sc_hd__decap_3 PHY_1067 ();
 sky130_fd_sc_hd__decap_3 PHY_1068 ();
 sky130_fd_sc_hd__decap_3 PHY_1069 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_1070 ();
 sky130_fd_sc_hd__decap_3 PHY_1071 ();
 sky130_fd_sc_hd__decap_3 PHY_1072 ();
 sky130_fd_sc_hd__decap_3 PHY_1073 ();
 sky130_fd_sc_hd__decap_3 PHY_1074 ();
 sky130_fd_sc_hd__decap_3 PHY_1075 ();
 sky130_fd_sc_hd__decap_3 PHY_1076 ();
 sky130_fd_sc_hd__decap_3 PHY_1077 ();
 sky130_fd_sc_hd__decap_3 PHY_1078 ();
 sky130_fd_sc_hd__decap_3 PHY_1079 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_1080 ();
 sky130_fd_sc_hd__decap_3 PHY_1081 ();
 sky130_fd_sc_hd__decap_3 PHY_1082 ();
 sky130_fd_sc_hd__decap_3 PHY_1083 ();
 sky130_fd_sc_hd__decap_3 PHY_1084 ();
 sky130_fd_sc_hd__decap_3 PHY_1085 ();
 sky130_fd_sc_hd__decap_3 PHY_1086 ();
 sky130_fd_sc_hd__decap_3 PHY_1087 ();
 sky130_fd_sc_hd__decap_3 PHY_1088 ();
 sky130_fd_sc_hd__decap_3 PHY_1089 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_1090 ();
 sky130_fd_sc_hd__decap_3 PHY_1091 ();
 sky130_fd_sc_hd__decap_3 PHY_1092 ();
 sky130_fd_sc_hd__decap_3 PHY_1093 ();
 sky130_fd_sc_hd__decap_3 PHY_1094 ();
 sky130_fd_sc_hd__decap_3 PHY_1095 ();
 sky130_fd_sc_hd__decap_3 PHY_1096 ();
 sky130_fd_sc_hd__decap_3 PHY_1097 ();
 sky130_fd_sc_hd__decap_3 PHY_1098 ();
 sky130_fd_sc_hd__decap_3 PHY_1099 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_1100 ();
 sky130_fd_sc_hd__decap_3 PHY_1101 ();
 sky130_fd_sc_hd__decap_3 PHY_1102 ();
 sky130_fd_sc_hd__decap_3 PHY_1103 ();
 sky130_fd_sc_hd__decap_3 PHY_1104 ();
 sky130_fd_sc_hd__decap_3 PHY_1105 ();
 sky130_fd_sc_hd__decap_3 PHY_1106 ();
 sky130_fd_sc_hd__decap_3 PHY_1107 ();
 sky130_fd_sc_hd__decap_3 PHY_1108 ();
 sky130_fd_sc_hd__decap_3 PHY_1109 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_1110 ();
 sky130_fd_sc_hd__decap_3 PHY_1111 ();
 sky130_fd_sc_hd__decap_3 PHY_1112 ();
 sky130_fd_sc_hd__decap_3 PHY_1113 ();
 sky130_fd_sc_hd__decap_3 PHY_1114 ();
 sky130_fd_sc_hd__decap_3 PHY_1115 ();
 sky130_fd_sc_hd__decap_3 PHY_1116 ();
 sky130_fd_sc_hd__decap_3 PHY_1117 ();
 sky130_fd_sc_hd__decap_3 PHY_1118 ();
 sky130_fd_sc_hd__decap_3 PHY_1119 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_1120 ();
 sky130_fd_sc_hd__decap_3 PHY_1121 ();
 sky130_fd_sc_hd__decap_3 PHY_1122 ();
 sky130_fd_sc_hd__decap_3 PHY_1123 ();
 sky130_fd_sc_hd__decap_3 PHY_1124 ();
 sky130_fd_sc_hd__decap_3 PHY_1125 ();
 sky130_fd_sc_hd__decap_3 PHY_1126 ();
 sky130_fd_sc_hd__decap_3 PHY_1127 ();
 sky130_fd_sc_hd__decap_3 PHY_1128 ();
 sky130_fd_sc_hd__decap_3 PHY_1129 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_1130 ();
 sky130_fd_sc_hd__decap_3 PHY_1131 ();
 sky130_fd_sc_hd__decap_3 PHY_1132 ();
 sky130_fd_sc_hd__decap_3 PHY_1133 ();
 sky130_fd_sc_hd__decap_3 PHY_1134 ();
 sky130_fd_sc_hd__decap_3 PHY_1135 ();
 sky130_fd_sc_hd__decap_3 PHY_1136 ();
 sky130_fd_sc_hd__decap_3 PHY_1137 ();
 sky130_fd_sc_hd__decap_3 PHY_1138 ();
 sky130_fd_sc_hd__decap_3 PHY_1139 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_1140 ();
 sky130_fd_sc_hd__decap_3 PHY_1141 ();
 sky130_fd_sc_hd__decap_3 PHY_1142 ();
 sky130_fd_sc_hd__decap_3 PHY_1143 ();
 sky130_fd_sc_hd__decap_3 PHY_1144 ();
 sky130_fd_sc_hd__decap_3 PHY_1145 ();
 sky130_fd_sc_hd__decap_3 PHY_1146 ();
 sky130_fd_sc_hd__decap_3 PHY_1147 ();
 sky130_fd_sc_hd__decap_3 PHY_1148 ();
 sky130_fd_sc_hd__decap_3 PHY_1149 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_1150 ();
 sky130_fd_sc_hd__decap_3 PHY_1151 ();
 sky130_fd_sc_hd__decap_3 PHY_1152 ();
 sky130_fd_sc_hd__decap_3 PHY_1153 ();
 sky130_fd_sc_hd__decap_3 PHY_1154 ();
 sky130_fd_sc_hd__decap_3 PHY_1155 ();
 sky130_fd_sc_hd__decap_3 PHY_1156 ();
 sky130_fd_sc_hd__decap_3 PHY_1157 ();
 sky130_fd_sc_hd__decap_3 PHY_1158 ();
 sky130_fd_sc_hd__decap_3 PHY_1159 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_1160 ();
 sky130_fd_sc_hd__decap_3 PHY_1161 ();
 sky130_fd_sc_hd__decap_3 PHY_1162 ();
 sky130_fd_sc_hd__decap_3 PHY_1163 ();
 sky130_fd_sc_hd__decap_3 PHY_1164 ();
 sky130_fd_sc_hd__decap_3 PHY_1165 ();
 sky130_fd_sc_hd__decap_3 PHY_1166 ();
 sky130_fd_sc_hd__decap_3 PHY_1167 ();
 sky130_fd_sc_hd__decap_3 PHY_1168 ();
 sky130_fd_sc_hd__decap_3 PHY_1169 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_1170 ();
 sky130_fd_sc_hd__decap_3 PHY_1171 ();
 sky130_fd_sc_hd__decap_3 PHY_1172 ();
 sky130_fd_sc_hd__decap_3 PHY_1173 ();
 sky130_fd_sc_hd__decap_3 PHY_1174 ();
 sky130_fd_sc_hd__decap_3 PHY_1175 ();
 sky130_fd_sc_hd__decap_3 PHY_1176 ();
 sky130_fd_sc_hd__decap_3 PHY_1177 ();
 sky130_fd_sc_hd__decap_3 PHY_1178 ();
 sky130_fd_sc_hd__decap_3 PHY_1179 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_1180 ();
 sky130_fd_sc_hd__decap_3 PHY_1181 ();
 sky130_fd_sc_hd__decap_3 PHY_1182 ();
 sky130_fd_sc_hd__decap_3 PHY_1183 ();
 sky130_fd_sc_hd__decap_3 PHY_1184 ();
 sky130_fd_sc_hd__decap_3 PHY_1185 ();
 sky130_fd_sc_hd__decap_3 PHY_1186 ();
 sky130_fd_sc_hd__decap_3 PHY_1187 ();
 sky130_fd_sc_hd__decap_3 PHY_1188 ();
 sky130_fd_sc_hd__decap_3 PHY_1189 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_1190 ();
 sky130_fd_sc_hd__decap_3 PHY_1191 ();
 sky130_fd_sc_hd__decap_3 PHY_1192 ();
 sky130_fd_sc_hd__decap_3 PHY_1193 ();
 sky130_fd_sc_hd__decap_3 PHY_1194 ();
 sky130_fd_sc_hd__decap_3 PHY_1195 ();
 sky130_fd_sc_hd__decap_3 PHY_1196 ();
 sky130_fd_sc_hd__decap_3 PHY_1197 ();
 sky130_fd_sc_hd__decap_3 PHY_1198 ();
 sky130_fd_sc_hd__decap_3 PHY_1199 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_1200 ();
 sky130_fd_sc_hd__decap_3 PHY_1201 ();
 sky130_fd_sc_hd__decap_3 PHY_1202 ();
 sky130_fd_sc_hd__decap_3 PHY_1203 ();
 sky130_fd_sc_hd__decap_3 PHY_1204 ();
 sky130_fd_sc_hd__decap_3 PHY_1205 ();
 sky130_fd_sc_hd__decap_3 PHY_1206 ();
 sky130_fd_sc_hd__decap_3 PHY_1207 ();
 sky130_fd_sc_hd__decap_3 PHY_1208 ();
 sky130_fd_sc_hd__decap_3 PHY_1209 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_1210 ();
 sky130_fd_sc_hd__decap_3 PHY_1211 ();
 sky130_fd_sc_hd__decap_3 PHY_1212 ();
 sky130_fd_sc_hd__decap_3 PHY_1213 ();
 sky130_fd_sc_hd__decap_3 PHY_1214 ();
 sky130_fd_sc_hd__decap_3 PHY_1215 ();
 sky130_fd_sc_hd__decap_3 PHY_1216 ();
 sky130_fd_sc_hd__decap_3 PHY_1217 ();
 sky130_fd_sc_hd__decap_3 PHY_1218 ();
 sky130_fd_sc_hd__decap_3 PHY_1219 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_1220 ();
 sky130_fd_sc_hd__decap_3 PHY_1221 ();
 sky130_fd_sc_hd__decap_3 PHY_1222 ();
 sky130_fd_sc_hd__decap_3 PHY_1223 ();
 sky130_fd_sc_hd__decap_3 PHY_1224 ();
 sky130_fd_sc_hd__decap_3 PHY_1225 ();
 sky130_fd_sc_hd__decap_3 PHY_1226 ();
 sky130_fd_sc_hd__decap_3 PHY_1227 ();
 sky130_fd_sc_hd__decap_3 PHY_1228 ();
 sky130_fd_sc_hd__decap_3 PHY_1229 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_1230 ();
 sky130_fd_sc_hd__decap_3 PHY_1231 ();
 sky130_fd_sc_hd__decap_3 PHY_1232 ();
 sky130_fd_sc_hd__decap_3 PHY_1233 ();
 sky130_fd_sc_hd__decap_3 PHY_1234 ();
 sky130_fd_sc_hd__decap_3 PHY_1235 ();
 sky130_fd_sc_hd__decap_3 PHY_1236 ();
 sky130_fd_sc_hd__decap_3 PHY_1237 ();
 sky130_fd_sc_hd__decap_3 PHY_1238 ();
 sky130_fd_sc_hd__decap_3 PHY_1239 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_1240 ();
 sky130_fd_sc_hd__decap_3 PHY_1241 ();
 sky130_fd_sc_hd__decap_3 PHY_1242 ();
 sky130_fd_sc_hd__decap_3 PHY_1243 ();
 sky130_fd_sc_hd__decap_3 PHY_1244 ();
 sky130_fd_sc_hd__decap_3 PHY_1245 ();
 sky130_fd_sc_hd__decap_3 PHY_1246 ();
 sky130_fd_sc_hd__decap_3 PHY_1247 ();
 sky130_fd_sc_hd__decap_3 PHY_1248 ();
 sky130_fd_sc_hd__decap_3 PHY_1249 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_1250 ();
 sky130_fd_sc_hd__decap_3 PHY_1251 ();
 sky130_fd_sc_hd__decap_3 PHY_1252 ();
 sky130_fd_sc_hd__decap_3 PHY_1253 ();
 sky130_fd_sc_hd__decap_3 PHY_1254 ();
 sky130_fd_sc_hd__decap_3 PHY_1255 ();
 sky130_fd_sc_hd__decap_3 PHY_1256 ();
 sky130_fd_sc_hd__decap_3 PHY_1257 ();
 sky130_fd_sc_hd__decap_3 PHY_1258 ();
 sky130_fd_sc_hd__decap_3 PHY_1259 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_1260 ();
 sky130_fd_sc_hd__decap_3 PHY_1261 ();
 sky130_fd_sc_hd__decap_3 PHY_1262 ();
 sky130_fd_sc_hd__decap_3 PHY_1263 ();
 sky130_fd_sc_hd__decap_3 PHY_1264 ();
 sky130_fd_sc_hd__decap_3 PHY_1265 ();
 sky130_fd_sc_hd__decap_3 PHY_1266 ();
 sky130_fd_sc_hd__decap_3 PHY_1267 ();
 sky130_fd_sc_hd__decap_3 PHY_1268 ();
 sky130_fd_sc_hd__decap_3 PHY_1269 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_1270 ();
 sky130_fd_sc_hd__decap_3 PHY_1271 ();
 sky130_fd_sc_hd__decap_3 PHY_1272 ();
 sky130_fd_sc_hd__decap_3 PHY_1273 ();
 sky130_fd_sc_hd__decap_3 PHY_1274 ();
 sky130_fd_sc_hd__decap_3 PHY_1275 ();
 sky130_fd_sc_hd__decap_3 PHY_1276 ();
 sky130_fd_sc_hd__decap_3 PHY_1277 ();
 sky130_fd_sc_hd__decap_3 PHY_1278 ();
 sky130_fd_sc_hd__decap_3 PHY_1279 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_1280 ();
 sky130_fd_sc_hd__decap_3 PHY_1281 ();
 sky130_fd_sc_hd__decap_3 PHY_1282 ();
 sky130_fd_sc_hd__decap_3 PHY_1283 ();
 sky130_fd_sc_hd__decap_3 PHY_1284 ();
 sky130_fd_sc_hd__decap_3 PHY_1285 ();
 sky130_fd_sc_hd__decap_3 PHY_1286 ();
 sky130_fd_sc_hd__decap_3 PHY_1287 ();
 sky130_fd_sc_hd__decap_3 PHY_1288 ();
 sky130_fd_sc_hd__decap_3 PHY_1289 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_1290 ();
 sky130_fd_sc_hd__decap_3 PHY_1291 ();
 sky130_fd_sc_hd__decap_3 PHY_1292 ();
 sky130_fd_sc_hd__decap_3 PHY_1293 ();
 sky130_fd_sc_hd__decap_3 PHY_1294 ();
 sky130_fd_sc_hd__decap_3 PHY_1295 ();
 sky130_fd_sc_hd__decap_3 PHY_1296 ();
 sky130_fd_sc_hd__decap_3 PHY_1297 ();
 sky130_fd_sc_hd__decap_3 PHY_1298 ();
 sky130_fd_sc_hd__decap_3 PHY_1299 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_1300 ();
 sky130_fd_sc_hd__decap_3 PHY_1301 ();
 sky130_fd_sc_hd__decap_3 PHY_1302 ();
 sky130_fd_sc_hd__decap_3 PHY_1303 ();
 sky130_fd_sc_hd__decap_3 PHY_1304 ();
 sky130_fd_sc_hd__decap_3 PHY_1305 ();
 sky130_fd_sc_hd__decap_3 PHY_1306 ();
 sky130_fd_sc_hd__decap_3 PHY_1307 ();
 sky130_fd_sc_hd__decap_3 PHY_1308 ();
 sky130_fd_sc_hd__decap_3 PHY_1309 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_1310 ();
 sky130_fd_sc_hd__decap_3 PHY_1311 ();
 sky130_fd_sc_hd__decap_3 PHY_1312 ();
 sky130_fd_sc_hd__decap_3 PHY_1313 ();
 sky130_fd_sc_hd__decap_3 PHY_1314 ();
 sky130_fd_sc_hd__decap_3 PHY_1315 ();
 sky130_fd_sc_hd__decap_3 PHY_1316 ();
 sky130_fd_sc_hd__decap_3 PHY_1317 ();
 sky130_fd_sc_hd__decap_3 PHY_1318 ();
 sky130_fd_sc_hd__decap_3 PHY_1319 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_1320 ();
 sky130_fd_sc_hd__decap_3 PHY_1321 ();
 sky130_fd_sc_hd__decap_3 PHY_1322 ();
 sky130_fd_sc_hd__decap_3 PHY_1323 ();
 sky130_fd_sc_hd__decap_3 PHY_1324 ();
 sky130_fd_sc_hd__decap_3 PHY_1325 ();
 sky130_fd_sc_hd__decap_3 PHY_1326 ();
 sky130_fd_sc_hd__decap_3 PHY_1327 ();
 sky130_fd_sc_hd__decap_3 PHY_1328 ();
 sky130_fd_sc_hd__decap_3 PHY_1329 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_1330 ();
 sky130_fd_sc_hd__decap_3 PHY_1331 ();
 sky130_fd_sc_hd__decap_3 PHY_1332 ();
 sky130_fd_sc_hd__decap_3 PHY_1333 ();
 sky130_fd_sc_hd__decap_3 PHY_1334 ();
 sky130_fd_sc_hd__decap_3 PHY_1335 ();
 sky130_fd_sc_hd__decap_3 PHY_1336 ();
 sky130_fd_sc_hd__decap_3 PHY_1337 ();
 sky130_fd_sc_hd__decap_3 PHY_1338 ();
 sky130_fd_sc_hd__decap_3 PHY_1339 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_1340 ();
 sky130_fd_sc_hd__decap_3 PHY_1341 ();
 sky130_fd_sc_hd__decap_3 PHY_1342 ();
 sky130_fd_sc_hd__decap_3 PHY_1343 ();
 sky130_fd_sc_hd__decap_3 PHY_1344 ();
 sky130_fd_sc_hd__decap_3 PHY_1345 ();
 sky130_fd_sc_hd__decap_3 PHY_1346 ();
 sky130_fd_sc_hd__decap_3 PHY_1347 ();
 sky130_fd_sc_hd__decap_3 PHY_1348 ();
 sky130_fd_sc_hd__decap_3 PHY_1349 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_1350 ();
 sky130_fd_sc_hd__decap_3 PHY_1351 ();
 sky130_fd_sc_hd__decap_3 PHY_1352 ();
 sky130_fd_sc_hd__decap_3 PHY_1353 ();
 sky130_fd_sc_hd__decap_3 PHY_1354 ();
 sky130_fd_sc_hd__decap_3 PHY_1355 ();
 sky130_fd_sc_hd__decap_3 PHY_1356 ();
 sky130_fd_sc_hd__decap_3 PHY_1357 ();
 sky130_fd_sc_hd__decap_3 PHY_1358 ();
 sky130_fd_sc_hd__decap_3 PHY_1359 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_1360 ();
 sky130_fd_sc_hd__decap_3 PHY_1361 ();
 sky130_fd_sc_hd__decap_3 PHY_1362 ();
 sky130_fd_sc_hd__decap_3 PHY_1363 ();
 sky130_fd_sc_hd__decap_3 PHY_1364 ();
 sky130_fd_sc_hd__decap_3 PHY_1365 ();
 sky130_fd_sc_hd__decap_3 PHY_1366 ();
 sky130_fd_sc_hd__decap_3 PHY_1367 ();
 sky130_fd_sc_hd__decap_3 PHY_1368 ();
 sky130_fd_sc_hd__decap_3 PHY_1369 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_1370 ();
 sky130_fd_sc_hd__decap_3 PHY_1371 ();
 sky130_fd_sc_hd__decap_3 PHY_1372 ();
 sky130_fd_sc_hd__decap_3 PHY_1373 ();
 sky130_fd_sc_hd__decap_3 PHY_1374 ();
 sky130_fd_sc_hd__decap_3 PHY_1375 ();
 sky130_fd_sc_hd__decap_3 PHY_1376 ();
 sky130_fd_sc_hd__decap_3 PHY_1377 ();
 sky130_fd_sc_hd__decap_3 PHY_1378 ();
 sky130_fd_sc_hd__decap_3 PHY_1379 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_1380 ();
 sky130_fd_sc_hd__decap_3 PHY_1381 ();
 sky130_fd_sc_hd__decap_3 PHY_1382 ();
 sky130_fd_sc_hd__decap_3 PHY_1383 ();
 sky130_fd_sc_hd__decap_3 PHY_1384 ();
 sky130_fd_sc_hd__decap_3 PHY_1385 ();
 sky130_fd_sc_hd__decap_3 PHY_1386 ();
 sky130_fd_sc_hd__decap_3 PHY_1387 ();
 sky130_fd_sc_hd__decap_3 PHY_1388 ();
 sky130_fd_sc_hd__decap_3 PHY_1389 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_1390 ();
 sky130_fd_sc_hd__decap_3 PHY_1391 ();
 sky130_fd_sc_hd__decap_3 PHY_1392 ();
 sky130_fd_sc_hd__decap_3 PHY_1393 ();
 sky130_fd_sc_hd__decap_3 PHY_1394 ();
 sky130_fd_sc_hd__decap_3 PHY_1395 ();
 sky130_fd_sc_hd__decap_3 PHY_1396 ();
 sky130_fd_sc_hd__decap_3 PHY_1397 ();
 sky130_fd_sc_hd__decap_3 PHY_1398 ();
 sky130_fd_sc_hd__decap_3 PHY_1399 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_1400 ();
 sky130_fd_sc_hd__decap_3 PHY_1401 ();
 sky130_fd_sc_hd__decap_3 PHY_1402 ();
 sky130_fd_sc_hd__decap_3 PHY_1403 ();
 sky130_fd_sc_hd__decap_3 PHY_1404 ();
 sky130_fd_sc_hd__decap_3 PHY_1405 ();
 sky130_fd_sc_hd__decap_3 PHY_1406 ();
 sky130_fd_sc_hd__decap_3 PHY_1407 ();
 sky130_fd_sc_hd__decap_3 PHY_1408 ();
 sky130_fd_sc_hd__decap_3 PHY_1409 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_1410 ();
 sky130_fd_sc_hd__decap_3 PHY_1411 ();
 sky130_fd_sc_hd__decap_3 PHY_1412 ();
 sky130_fd_sc_hd__decap_3 PHY_1413 ();
 sky130_fd_sc_hd__decap_3 PHY_1414 ();
 sky130_fd_sc_hd__decap_3 PHY_1415 ();
 sky130_fd_sc_hd__decap_3 PHY_1416 ();
 sky130_fd_sc_hd__decap_3 PHY_1417 ();
 sky130_fd_sc_hd__decap_3 PHY_1418 ();
 sky130_fd_sc_hd__decap_3 PHY_1419 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_1420 ();
 sky130_fd_sc_hd__decap_3 PHY_1421 ();
 sky130_fd_sc_hd__decap_3 PHY_1422 ();
 sky130_fd_sc_hd__decap_3 PHY_1423 ();
 sky130_fd_sc_hd__decap_3 PHY_1424 ();
 sky130_fd_sc_hd__decap_3 PHY_1425 ();
 sky130_fd_sc_hd__decap_3 PHY_1426 ();
 sky130_fd_sc_hd__decap_3 PHY_1427 ();
 sky130_fd_sc_hd__decap_3 PHY_1428 ();
 sky130_fd_sc_hd__decap_3 PHY_1429 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_1430 ();
 sky130_fd_sc_hd__decap_3 PHY_1431 ();
 sky130_fd_sc_hd__decap_3 PHY_1432 ();
 sky130_fd_sc_hd__decap_3 PHY_1433 ();
 sky130_fd_sc_hd__decap_3 PHY_1434 ();
 sky130_fd_sc_hd__decap_3 PHY_1435 ();
 sky130_fd_sc_hd__decap_3 PHY_1436 ();
 sky130_fd_sc_hd__decap_3 PHY_1437 ();
 sky130_fd_sc_hd__decap_3 PHY_1438 ();
 sky130_fd_sc_hd__decap_3 PHY_1439 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_1440 ();
 sky130_fd_sc_hd__decap_3 PHY_1441 ();
 sky130_fd_sc_hd__decap_3 PHY_1442 ();
 sky130_fd_sc_hd__decap_3 PHY_1443 ();
 sky130_fd_sc_hd__decap_3 PHY_1444 ();
 sky130_fd_sc_hd__decap_3 PHY_1445 ();
 sky130_fd_sc_hd__decap_3 PHY_1446 ();
 sky130_fd_sc_hd__decap_3 PHY_1447 ();
 sky130_fd_sc_hd__decap_3 PHY_1448 ();
 sky130_fd_sc_hd__decap_3 PHY_1449 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_1450 ();
 sky130_fd_sc_hd__decap_3 PHY_1451 ();
 sky130_fd_sc_hd__decap_3 PHY_1452 ();
 sky130_fd_sc_hd__decap_3 PHY_1453 ();
 sky130_fd_sc_hd__decap_3 PHY_1454 ();
 sky130_fd_sc_hd__decap_3 PHY_1455 ();
 sky130_fd_sc_hd__decap_3 PHY_1456 ();
 sky130_fd_sc_hd__decap_3 PHY_1457 ();
 sky130_fd_sc_hd__decap_3 PHY_1458 ();
 sky130_fd_sc_hd__decap_3 PHY_1459 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_1460 ();
 sky130_fd_sc_hd__decap_3 PHY_1461 ();
 sky130_fd_sc_hd__decap_3 PHY_1462 ();
 sky130_fd_sc_hd__decap_3 PHY_1463 ();
 sky130_fd_sc_hd__decap_3 PHY_1464 ();
 sky130_fd_sc_hd__decap_3 PHY_1465 ();
 sky130_fd_sc_hd__decap_3 PHY_1466 ();
 sky130_fd_sc_hd__decap_3 PHY_1467 ();
 sky130_fd_sc_hd__decap_3 PHY_1468 ();
 sky130_fd_sc_hd__decap_3 PHY_1469 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_1470 ();
 sky130_fd_sc_hd__decap_3 PHY_1471 ();
 sky130_fd_sc_hd__decap_3 PHY_1472 ();
 sky130_fd_sc_hd__decap_3 PHY_1473 ();
 sky130_fd_sc_hd__decap_3 PHY_1474 ();
 sky130_fd_sc_hd__decap_3 PHY_1475 ();
 sky130_fd_sc_hd__decap_3 PHY_1476 ();
 sky130_fd_sc_hd__decap_3 PHY_1477 ();
 sky130_fd_sc_hd__decap_3 PHY_1478 ();
 sky130_fd_sc_hd__decap_3 PHY_1479 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_1480 ();
 sky130_fd_sc_hd__decap_3 PHY_1481 ();
 sky130_fd_sc_hd__decap_3 PHY_1482 ();
 sky130_fd_sc_hd__decap_3 PHY_1483 ();
 sky130_fd_sc_hd__decap_3 PHY_1484 ();
 sky130_fd_sc_hd__decap_3 PHY_1485 ();
 sky130_fd_sc_hd__decap_3 PHY_1486 ();
 sky130_fd_sc_hd__decap_3 PHY_1487 ();
 sky130_fd_sc_hd__decap_3 PHY_1488 ();
 sky130_fd_sc_hd__decap_3 PHY_1489 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_1490 ();
 sky130_fd_sc_hd__decap_3 PHY_1491 ();
 sky130_fd_sc_hd__decap_3 PHY_1492 ();
 sky130_fd_sc_hd__decap_3 PHY_1493 ();
 sky130_fd_sc_hd__decap_3 PHY_1494 ();
 sky130_fd_sc_hd__decap_3 PHY_1495 ();
 sky130_fd_sc_hd__decap_3 PHY_1496 ();
 sky130_fd_sc_hd__decap_3 PHY_1497 ();
 sky130_fd_sc_hd__decap_3 PHY_1498 ();
 sky130_fd_sc_hd__decap_3 PHY_1499 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_1500 ();
 sky130_fd_sc_hd__decap_3 PHY_1501 ();
 sky130_fd_sc_hd__decap_3 PHY_1502 ();
 sky130_fd_sc_hd__decap_3 PHY_1503 ();
 sky130_fd_sc_hd__decap_3 PHY_1504 ();
 sky130_fd_sc_hd__decap_3 PHY_1505 ();
 sky130_fd_sc_hd__decap_3 PHY_1506 ();
 sky130_fd_sc_hd__decap_3 PHY_1507 ();
 sky130_fd_sc_hd__decap_3 PHY_1508 ();
 sky130_fd_sc_hd__decap_3 PHY_1509 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_1510 ();
 sky130_fd_sc_hd__decap_3 PHY_1511 ();
 sky130_fd_sc_hd__decap_3 PHY_1512 ();
 sky130_fd_sc_hd__decap_3 PHY_1513 ();
 sky130_fd_sc_hd__decap_3 PHY_1514 ();
 sky130_fd_sc_hd__decap_3 PHY_1515 ();
 sky130_fd_sc_hd__decap_3 PHY_1516 ();
 sky130_fd_sc_hd__decap_3 PHY_1517 ();
 sky130_fd_sc_hd__decap_3 PHY_1518 ();
 sky130_fd_sc_hd__decap_3 PHY_1519 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_1520 ();
 sky130_fd_sc_hd__decap_3 PHY_1521 ();
 sky130_fd_sc_hd__decap_3 PHY_1522 ();
 sky130_fd_sc_hd__decap_3 PHY_1523 ();
 sky130_fd_sc_hd__decap_3 PHY_1524 ();
 sky130_fd_sc_hd__decap_3 PHY_1525 ();
 sky130_fd_sc_hd__decap_3 PHY_1526 ();
 sky130_fd_sc_hd__decap_3 PHY_1527 ();
 sky130_fd_sc_hd__decap_3 PHY_1528 ();
 sky130_fd_sc_hd__decap_3 PHY_1529 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_1530 ();
 sky130_fd_sc_hd__decap_3 PHY_1531 ();
 sky130_fd_sc_hd__decap_3 PHY_1532 ();
 sky130_fd_sc_hd__decap_3 PHY_1533 ();
 sky130_fd_sc_hd__decap_3 PHY_1534 ();
 sky130_fd_sc_hd__decap_3 PHY_1535 ();
 sky130_fd_sc_hd__decap_3 PHY_1536 ();
 sky130_fd_sc_hd__decap_3 PHY_1537 ();
 sky130_fd_sc_hd__decap_3 PHY_1538 ();
 sky130_fd_sc_hd__decap_3 PHY_1539 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_1540 ();
 sky130_fd_sc_hd__decap_3 PHY_1541 ();
 sky130_fd_sc_hd__decap_3 PHY_1542 ();
 sky130_fd_sc_hd__decap_3 PHY_1543 ();
 sky130_fd_sc_hd__decap_3 PHY_1544 ();
 sky130_fd_sc_hd__decap_3 PHY_1545 ();
 sky130_fd_sc_hd__decap_3 PHY_1546 ();
 sky130_fd_sc_hd__decap_3 PHY_1547 ();
 sky130_fd_sc_hd__decap_3 PHY_1548 ();
 sky130_fd_sc_hd__decap_3 PHY_1549 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_1550 ();
 sky130_fd_sc_hd__decap_3 PHY_1551 ();
 sky130_fd_sc_hd__decap_3 PHY_1552 ();
 sky130_fd_sc_hd__decap_3 PHY_1553 ();
 sky130_fd_sc_hd__decap_3 PHY_1554 ();
 sky130_fd_sc_hd__decap_3 PHY_1555 ();
 sky130_fd_sc_hd__decap_3 PHY_1556 ();
 sky130_fd_sc_hd__decap_3 PHY_1557 ();
 sky130_fd_sc_hd__decap_3 PHY_1558 ();
 sky130_fd_sc_hd__decap_3 PHY_1559 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_1560 ();
 sky130_fd_sc_hd__decap_3 PHY_1561 ();
 sky130_fd_sc_hd__decap_3 PHY_1562 ();
 sky130_fd_sc_hd__decap_3 PHY_1563 ();
 sky130_fd_sc_hd__decap_3 PHY_1564 ();
 sky130_fd_sc_hd__decap_3 PHY_1565 ();
 sky130_fd_sc_hd__decap_3 PHY_1566 ();
 sky130_fd_sc_hd__decap_3 PHY_1567 ();
 sky130_fd_sc_hd__decap_3 PHY_1568 ();
 sky130_fd_sc_hd__decap_3 PHY_1569 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_1570 ();
 sky130_fd_sc_hd__decap_3 PHY_1571 ();
 sky130_fd_sc_hd__decap_3 PHY_1572 ();
 sky130_fd_sc_hd__decap_3 PHY_1573 ();
 sky130_fd_sc_hd__decap_3 PHY_1574 ();
 sky130_fd_sc_hd__decap_3 PHY_1575 ();
 sky130_fd_sc_hd__decap_3 PHY_1576 ();
 sky130_fd_sc_hd__decap_3 PHY_1577 ();
 sky130_fd_sc_hd__decap_3 PHY_1578 ();
 sky130_fd_sc_hd__decap_3 PHY_1579 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_1580 ();
 sky130_fd_sc_hd__decap_3 PHY_1581 ();
 sky130_fd_sc_hd__decap_3 PHY_1582 ();
 sky130_fd_sc_hd__decap_3 PHY_1583 ();
 sky130_fd_sc_hd__decap_3 PHY_1584 ();
 sky130_fd_sc_hd__decap_3 PHY_1585 ();
 sky130_fd_sc_hd__decap_3 PHY_1586 ();
 sky130_fd_sc_hd__decap_3 PHY_1587 ();
 sky130_fd_sc_hd__decap_3 PHY_1588 ();
 sky130_fd_sc_hd__decap_3 PHY_1589 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_1590 ();
 sky130_fd_sc_hd__decap_3 PHY_1591 ();
 sky130_fd_sc_hd__decap_3 PHY_1592 ();
 sky130_fd_sc_hd__decap_3 PHY_1593 ();
 sky130_fd_sc_hd__decap_3 PHY_1594 ();
 sky130_fd_sc_hd__decap_3 PHY_1595 ();
 sky130_fd_sc_hd__decap_3 PHY_1596 ();
 sky130_fd_sc_hd__decap_3 PHY_1597 ();
 sky130_fd_sc_hd__decap_3 PHY_1598 ();
 sky130_fd_sc_hd__decap_3 PHY_1599 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_1600 ();
 sky130_fd_sc_hd__decap_3 PHY_1601 ();
 sky130_fd_sc_hd__decap_3 PHY_1602 ();
 sky130_fd_sc_hd__decap_3 PHY_1603 ();
 sky130_fd_sc_hd__decap_3 PHY_1604 ();
 sky130_fd_sc_hd__decap_3 PHY_1605 ();
 sky130_fd_sc_hd__decap_3 PHY_1606 ();
 sky130_fd_sc_hd__decap_3 PHY_1607 ();
 sky130_fd_sc_hd__decap_3 PHY_1608 ();
 sky130_fd_sc_hd__decap_3 PHY_1609 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_1610 ();
 sky130_fd_sc_hd__decap_3 PHY_1611 ();
 sky130_fd_sc_hd__decap_3 PHY_1612 ();
 sky130_fd_sc_hd__decap_3 PHY_1613 ();
 sky130_fd_sc_hd__decap_3 PHY_1614 ();
 sky130_fd_sc_hd__decap_3 PHY_1615 ();
 sky130_fd_sc_hd__decap_3 PHY_1616 ();
 sky130_fd_sc_hd__decap_3 PHY_1617 ();
 sky130_fd_sc_hd__decap_3 PHY_1618 ();
 sky130_fd_sc_hd__decap_3 PHY_1619 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_1620 ();
 sky130_fd_sc_hd__decap_3 PHY_1621 ();
 sky130_fd_sc_hd__decap_3 PHY_1622 ();
 sky130_fd_sc_hd__decap_3 PHY_1623 ();
 sky130_fd_sc_hd__decap_3 PHY_1624 ();
 sky130_fd_sc_hd__decap_3 PHY_1625 ();
 sky130_fd_sc_hd__decap_3 PHY_1626 ();
 sky130_fd_sc_hd__decap_3 PHY_1627 ();
 sky130_fd_sc_hd__decap_3 PHY_1628 ();
 sky130_fd_sc_hd__decap_3 PHY_1629 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_1630 ();
 sky130_fd_sc_hd__decap_3 PHY_1631 ();
 sky130_fd_sc_hd__decap_3 PHY_1632 ();
 sky130_fd_sc_hd__decap_3 PHY_1633 ();
 sky130_fd_sc_hd__decap_3 PHY_1634 ();
 sky130_fd_sc_hd__decap_3 PHY_1635 ();
 sky130_fd_sc_hd__decap_3 PHY_1636 ();
 sky130_fd_sc_hd__decap_3 PHY_1637 ();
 sky130_fd_sc_hd__decap_3 PHY_1638 ();
 sky130_fd_sc_hd__decap_3 PHY_1639 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_1640 ();
 sky130_fd_sc_hd__decap_3 PHY_1641 ();
 sky130_fd_sc_hd__decap_3 PHY_1642 ();
 sky130_fd_sc_hd__decap_3 PHY_1643 ();
 sky130_fd_sc_hd__decap_3 PHY_1644 ();
 sky130_fd_sc_hd__decap_3 PHY_1645 ();
 sky130_fd_sc_hd__decap_3 PHY_1646 ();
 sky130_fd_sc_hd__decap_3 PHY_1647 ();
 sky130_fd_sc_hd__decap_3 PHY_1648 ();
 sky130_fd_sc_hd__decap_3 PHY_1649 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_1650 ();
 sky130_fd_sc_hd__decap_3 PHY_1651 ();
 sky130_fd_sc_hd__decap_3 PHY_1652 ();
 sky130_fd_sc_hd__decap_3 PHY_1653 ();
 sky130_fd_sc_hd__decap_3 PHY_1654 ();
 sky130_fd_sc_hd__decap_3 PHY_1655 ();
 sky130_fd_sc_hd__decap_3 PHY_1656 ();
 sky130_fd_sc_hd__decap_3 PHY_1657 ();
 sky130_fd_sc_hd__decap_3 PHY_1658 ();
 sky130_fd_sc_hd__decap_3 PHY_1659 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_1660 ();
 sky130_fd_sc_hd__decap_3 PHY_1661 ();
 sky130_fd_sc_hd__decap_3 PHY_1662 ();
 sky130_fd_sc_hd__decap_3 PHY_1663 ();
 sky130_fd_sc_hd__decap_3 PHY_1664 ();
 sky130_fd_sc_hd__decap_3 PHY_1665 ();
 sky130_fd_sc_hd__decap_3 PHY_1666 ();
 sky130_fd_sc_hd__decap_3 PHY_1667 ();
 sky130_fd_sc_hd__decap_3 PHY_1668 ();
 sky130_fd_sc_hd__decap_3 PHY_1669 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_1670 ();
 sky130_fd_sc_hd__decap_3 PHY_1671 ();
 sky130_fd_sc_hd__decap_3 PHY_1672 ();
 sky130_fd_sc_hd__decap_3 PHY_1673 ();
 sky130_fd_sc_hd__decap_3 PHY_1674 ();
 sky130_fd_sc_hd__decap_3 PHY_1675 ();
 sky130_fd_sc_hd__decap_3 PHY_1676 ();
 sky130_fd_sc_hd__decap_3 PHY_1677 ();
 sky130_fd_sc_hd__decap_3 PHY_1678 ();
 sky130_fd_sc_hd__decap_3 PHY_1679 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_1680 ();
 sky130_fd_sc_hd__decap_3 PHY_1681 ();
 sky130_fd_sc_hd__decap_3 PHY_1682 ();
 sky130_fd_sc_hd__decap_3 PHY_1683 ();
 sky130_fd_sc_hd__decap_3 PHY_1684 ();
 sky130_fd_sc_hd__decap_3 PHY_1685 ();
 sky130_fd_sc_hd__decap_3 PHY_1686 ();
 sky130_fd_sc_hd__decap_3 PHY_1687 ();
 sky130_fd_sc_hd__decap_3 PHY_1688 ();
 sky130_fd_sc_hd__decap_3 PHY_1689 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_1690 ();
 sky130_fd_sc_hd__decap_3 PHY_1691 ();
 sky130_fd_sc_hd__decap_3 PHY_1692 ();
 sky130_fd_sc_hd__decap_3 PHY_1693 ();
 sky130_fd_sc_hd__decap_3 PHY_1694 ();
 sky130_fd_sc_hd__decap_3 PHY_1695 ();
 sky130_fd_sc_hd__decap_3 PHY_1696 ();
 sky130_fd_sc_hd__decap_3 PHY_1697 ();
 sky130_fd_sc_hd__decap_3 PHY_1698 ();
 sky130_fd_sc_hd__decap_3 PHY_1699 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_1700 ();
 sky130_fd_sc_hd__decap_3 PHY_1701 ();
 sky130_fd_sc_hd__decap_3 PHY_1702 ();
 sky130_fd_sc_hd__decap_3 PHY_1703 ();
 sky130_fd_sc_hd__decap_3 PHY_1704 ();
 sky130_fd_sc_hd__decap_3 PHY_1705 ();
 sky130_fd_sc_hd__decap_3 PHY_1706 ();
 sky130_fd_sc_hd__decap_3 PHY_1707 ();
 sky130_fd_sc_hd__decap_3 PHY_1708 ();
 sky130_fd_sc_hd__decap_3 PHY_1709 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_1710 ();
 sky130_fd_sc_hd__decap_3 PHY_1711 ();
 sky130_fd_sc_hd__decap_3 PHY_1712 ();
 sky130_fd_sc_hd__decap_3 PHY_1713 ();
 sky130_fd_sc_hd__decap_3 PHY_1714 ();
 sky130_fd_sc_hd__decap_3 PHY_1715 ();
 sky130_fd_sc_hd__decap_3 PHY_1716 ();
 sky130_fd_sc_hd__decap_3 PHY_1717 ();
 sky130_fd_sc_hd__decap_3 PHY_1718 ();
 sky130_fd_sc_hd__decap_3 PHY_1719 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_1720 ();
 sky130_fd_sc_hd__decap_3 PHY_1721 ();
 sky130_fd_sc_hd__decap_3 PHY_1722 ();
 sky130_fd_sc_hd__decap_3 PHY_1723 ();
 sky130_fd_sc_hd__decap_3 PHY_1724 ();
 sky130_fd_sc_hd__decap_3 PHY_1725 ();
 sky130_fd_sc_hd__decap_3 PHY_1726 ();
 sky130_fd_sc_hd__decap_3 PHY_1727 ();
 sky130_fd_sc_hd__decap_3 PHY_1728 ();
 sky130_fd_sc_hd__decap_3 PHY_1729 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_1730 ();
 sky130_fd_sc_hd__decap_3 PHY_1731 ();
 sky130_fd_sc_hd__decap_3 PHY_1732 ();
 sky130_fd_sc_hd__decap_3 PHY_1733 ();
 sky130_fd_sc_hd__decap_3 PHY_1734 ();
 sky130_fd_sc_hd__decap_3 PHY_1735 ();
 sky130_fd_sc_hd__decap_3 PHY_1736 ();
 sky130_fd_sc_hd__decap_3 PHY_1737 ();
 sky130_fd_sc_hd__decap_3 PHY_1738 ();
 sky130_fd_sc_hd__decap_3 PHY_1739 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_1740 ();
 sky130_fd_sc_hd__decap_3 PHY_1741 ();
 sky130_fd_sc_hd__decap_3 PHY_1742 ();
 sky130_fd_sc_hd__decap_3 PHY_1743 ();
 sky130_fd_sc_hd__decap_3 PHY_1744 ();
 sky130_fd_sc_hd__decap_3 PHY_1745 ();
 sky130_fd_sc_hd__decap_3 PHY_1746 ();
 sky130_fd_sc_hd__decap_3 PHY_1747 ();
 sky130_fd_sc_hd__decap_3 PHY_1748 ();
 sky130_fd_sc_hd__decap_3 PHY_1749 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_1750 ();
 sky130_fd_sc_hd__decap_3 PHY_1751 ();
 sky130_fd_sc_hd__decap_3 PHY_1752 ();
 sky130_fd_sc_hd__decap_3 PHY_1753 ();
 sky130_fd_sc_hd__decap_3 PHY_1754 ();
 sky130_fd_sc_hd__decap_3 PHY_1755 ();
 sky130_fd_sc_hd__decap_3 PHY_1756 ();
 sky130_fd_sc_hd__decap_3 PHY_1757 ();
 sky130_fd_sc_hd__decap_3 PHY_1758 ();
 sky130_fd_sc_hd__decap_3 PHY_1759 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_1760 ();
 sky130_fd_sc_hd__decap_3 PHY_1761 ();
 sky130_fd_sc_hd__decap_3 PHY_1762 ();
 sky130_fd_sc_hd__decap_3 PHY_1763 ();
 sky130_fd_sc_hd__decap_3 PHY_1764 ();
 sky130_fd_sc_hd__decap_3 PHY_1765 ();
 sky130_fd_sc_hd__decap_3 PHY_1766 ();
 sky130_fd_sc_hd__decap_3 PHY_1767 ();
 sky130_fd_sc_hd__decap_3 PHY_1768 ();
 sky130_fd_sc_hd__decap_3 PHY_1769 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_1770 ();
 sky130_fd_sc_hd__decap_3 PHY_1771 ();
 sky130_fd_sc_hd__decap_3 PHY_1772 ();
 sky130_fd_sc_hd__decap_3 PHY_1773 ();
 sky130_fd_sc_hd__decap_3 PHY_1774 ();
 sky130_fd_sc_hd__decap_3 PHY_1775 ();
 sky130_fd_sc_hd__decap_3 PHY_1776 ();
 sky130_fd_sc_hd__decap_3 PHY_1777 ();
 sky130_fd_sc_hd__decap_3 PHY_1778 ();
 sky130_fd_sc_hd__decap_3 PHY_1779 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_1780 ();
 sky130_fd_sc_hd__decap_3 PHY_1781 ();
 sky130_fd_sc_hd__decap_3 PHY_1782 ();
 sky130_fd_sc_hd__decap_3 PHY_1783 ();
 sky130_fd_sc_hd__decap_3 PHY_1784 ();
 sky130_fd_sc_hd__decap_3 PHY_1785 ();
 sky130_fd_sc_hd__decap_3 PHY_1786 ();
 sky130_fd_sc_hd__decap_3 PHY_1787 ();
 sky130_fd_sc_hd__decap_3 PHY_1788 ();
 sky130_fd_sc_hd__decap_3 PHY_1789 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_1790 ();
 sky130_fd_sc_hd__decap_3 PHY_1791 ();
 sky130_fd_sc_hd__decap_3 PHY_1792 ();
 sky130_fd_sc_hd__decap_3 PHY_1793 ();
 sky130_fd_sc_hd__decap_3 PHY_1794 ();
 sky130_fd_sc_hd__decap_3 PHY_1795 ();
 sky130_fd_sc_hd__decap_3 PHY_1796 ();
 sky130_fd_sc_hd__decap_3 PHY_1797 ();
 sky130_fd_sc_hd__decap_3 PHY_1798 ();
 sky130_fd_sc_hd__decap_3 PHY_1799 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_1800 ();
 sky130_fd_sc_hd__decap_3 PHY_1801 ();
 sky130_fd_sc_hd__decap_3 PHY_1802 ();
 sky130_fd_sc_hd__decap_3 PHY_1803 ();
 sky130_fd_sc_hd__decap_3 PHY_1804 ();
 sky130_fd_sc_hd__decap_3 PHY_1805 ();
 sky130_fd_sc_hd__decap_3 PHY_1806 ();
 sky130_fd_sc_hd__decap_3 PHY_1807 ();
 sky130_fd_sc_hd__decap_3 PHY_1808 ();
 sky130_fd_sc_hd__decap_3 PHY_1809 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_1810 ();
 sky130_fd_sc_hd__decap_3 PHY_1811 ();
 sky130_fd_sc_hd__decap_3 PHY_1812 ();
 sky130_fd_sc_hd__decap_3 PHY_1813 ();
 sky130_fd_sc_hd__decap_3 PHY_1814 ();
 sky130_fd_sc_hd__decap_3 PHY_1815 ();
 sky130_fd_sc_hd__decap_3 PHY_1816 ();
 sky130_fd_sc_hd__decap_3 PHY_1817 ();
 sky130_fd_sc_hd__decap_3 PHY_1818 ();
 sky130_fd_sc_hd__decap_3 PHY_1819 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_1820 ();
 sky130_fd_sc_hd__decap_3 PHY_1821 ();
 sky130_fd_sc_hd__decap_3 PHY_1822 ();
 sky130_fd_sc_hd__decap_3 PHY_1823 ();
 sky130_fd_sc_hd__decap_3 PHY_1824 ();
 sky130_fd_sc_hd__decap_3 PHY_1825 ();
 sky130_fd_sc_hd__decap_3 PHY_1826 ();
 sky130_fd_sc_hd__decap_3 PHY_1827 ();
 sky130_fd_sc_hd__decap_3 PHY_1828 ();
 sky130_fd_sc_hd__decap_3 PHY_1829 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_1830 ();
 sky130_fd_sc_hd__decap_3 PHY_1831 ();
 sky130_fd_sc_hd__decap_3 PHY_1832 ();
 sky130_fd_sc_hd__decap_3 PHY_1833 ();
 sky130_fd_sc_hd__decap_3 PHY_1834 ();
 sky130_fd_sc_hd__decap_3 PHY_1835 ();
 sky130_fd_sc_hd__decap_3 PHY_1836 ();
 sky130_fd_sc_hd__decap_3 PHY_1837 ();
 sky130_fd_sc_hd__decap_3 PHY_1838 ();
 sky130_fd_sc_hd__decap_3 PHY_1839 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_1840 ();
 sky130_fd_sc_hd__decap_3 PHY_1841 ();
 sky130_fd_sc_hd__decap_3 PHY_1842 ();
 sky130_fd_sc_hd__decap_3 PHY_1843 ();
 sky130_fd_sc_hd__decap_3 PHY_1844 ();
 sky130_fd_sc_hd__decap_3 PHY_1845 ();
 sky130_fd_sc_hd__decap_3 PHY_1846 ();
 sky130_fd_sc_hd__decap_3 PHY_1847 ();
 sky130_fd_sc_hd__decap_3 PHY_1848 ();
 sky130_fd_sc_hd__decap_3 PHY_1849 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_1850 ();
 sky130_fd_sc_hd__decap_3 PHY_1851 ();
 sky130_fd_sc_hd__decap_3 PHY_1852 ();
 sky130_fd_sc_hd__decap_3 PHY_1853 ();
 sky130_fd_sc_hd__decap_3 PHY_1854 ();
 sky130_fd_sc_hd__decap_3 PHY_1855 ();
 sky130_fd_sc_hd__decap_3 PHY_1856 ();
 sky130_fd_sc_hd__decap_3 PHY_1857 ();
 sky130_fd_sc_hd__decap_3 PHY_1858 ();
 sky130_fd_sc_hd__decap_3 PHY_1859 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_1860 ();
 sky130_fd_sc_hd__decap_3 PHY_1861 ();
 sky130_fd_sc_hd__decap_3 PHY_1862 ();
 sky130_fd_sc_hd__decap_3 PHY_1863 ();
 sky130_fd_sc_hd__decap_3 PHY_1864 ();
 sky130_fd_sc_hd__decap_3 PHY_1865 ();
 sky130_fd_sc_hd__decap_3 PHY_1866 ();
 sky130_fd_sc_hd__decap_3 PHY_1867 ();
 sky130_fd_sc_hd__decap_3 PHY_1868 ();
 sky130_fd_sc_hd__decap_3 PHY_1869 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_1870 ();
 sky130_fd_sc_hd__decap_3 PHY_1871 ();
 sky130_fd_sc_hd__decap_3 PHY_1872 ();
 sky130_fd_sc_hd__decap_3 PHY_1873 ();
 sky130_fd_sc_hd__decap_3 PHY_1874 ();
 sky130_fd_sc_hd__decap_3 PHY_1875 ();
 sky130_fd_sc_hd__decap_3 PHY_1876 ();
 sky130_fd_sc_hd__decap_3 PHY_1877 ();
 sky130_fd_sc_hd__decap_3 PHY_1878 ();
 sky130_fd_sc_hd__decap_3 PHY_1879 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_1880 ();
 sky130_fd_sc_hd__decap_3 PHY_1881 ();
 sky130_fd_sc_hd__decap_3 PHY_1882 ();
 sky130_fd_sc_hd__decap_3 PHY_1883 ();
 sky130_fd_sc_hd__decap_3 PHY_1884 ();
 sky130_fd_sc_hd__decap_3 PHY_1885 ();
 sky130_fd_sc_hd__decap_3 PHY_1886 ();
 sky130_fd_sc_hd__decap_3 PHY_1887 ();
 sky130_fd_sc_hd__decap_3 PHY_1888 ();
 sky130_fd_sc_hd__decap_3 PHY_1889 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_1890 ();
 sky130_fd_sc_hd__decap_3 PHY_1891 ();
 sky130_fd_sc_hd__decap_3 PHY_1892 ();
 sky130_fd_sc_hd__decap_3 PHY_1893 ();
 sky130_fd_sc_hd__decap_3 PHY_1894 ();
 sky130_fd_sc_hd__decap_3 PHY_1895 ();
 sky130_fd_sc_hd__decap_3 PHY_1896 ();
 sky130_fd_sc_hd__decap_3 PHY_1897 ();
 sky130_fd_sc_hd__decap_3 PHY_1898 ();
 sky130_fd_sc_hd__decap_3 PHY_1899 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_1900 ();
 sky130_fd_sc_hd__decap_3 PHY_1901 ();
 sky130_fd_sc_hd__decap_3 PHY_1902 ();
 sky130_fd_sc_hd__decap_3 PHY_1903 ();
 sky130_fd_sc_hd__decap_3 PHY_1904 ();
 sky130_fd_sc_hd__decap_3 PHY_1905 ();
 sky130_fd_sc_hd__decap_3 PHY_1906 ();
 sky130_fd_sc_hd__decap_3 PHY_1907 ();
 sky130_fd_sc_hd__decap_3 PHY_1908 ();
 sky130_fd_sc_hd__decap_3 PHY_1909 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_1910 ();
 sky130_fd_sc_hd__decap_3 PHY_1911 ();
 sky130_fd_sc_hd__decap_3 PHY_1912 ();
 sky130_fd_sc_hd__decap_3 PHY_1913 ();
 sky130_fd_sc_hd__decap_3 PHY_1914 ();
 sky130_fd_sc_hd__decap_3 PHY_1915 ();
 sky130_fd_sc_hd__decap_3 PHY_1916 ();
 sky130_fd_sc_hd__decap_3 PHY_1917 ();
 sky130_fd_sc_hd__decap_3 PHY_1918 ();
 sky130_fd_sc_hd__decap_3 PHY_1919 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_1920 ();
 sky130_fd_sc_hd__decap_3 PHY_1921 ();
 sky130_fd_sc_hd__decap_3 PHY_1922 ();
 sky130_fd_sc_hd__decap_3 PHY_1923 ();
 sky130_fd_sc_hd__decap_3 PHY_1924 ();
 sky130_fd_sc_hd__decap_3 PHY_1925 ();
 sky130_fd_sc_hd__decap_3 PHY_1926 ();
 sky130_fd_sc_hd__decap_3 PHY_1927 ();
 sky130_fd_sc_hd__decap_3 PHY_1928 ();
 sky130_fd_sc_hd__decap_3 PHY_1929 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_1930 ();
 sky130_fd_sc_hd__decap_3 PHY_1931 ();
 sky130_fd_sc_hd__decap_3 PHY_1932 ();
 sky130_fd_sc_hd__decap_3 PHY_1933 ();
 sky130_fd_sc_hd__decap_3 PHY_1934 ();
 sky130_fd_sc_hd__decap_3 PHY_1935 ();
 sky130_fd_sc_hd__decap_3 PHY_1936 ();
 sky130_fd_sc_hd__decap_3 PHY_1937 ();
 sky130_fd_sc_hd__decap_3 PHY_1938 ();
 sky130_fd_sc_hd__decap_3 PHY_1939 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_1940 ();
 sky130_fd_sc_hd__decap_3 PHY_1941 ();
 sky130_fd_sc_hd__decap_3 PHY_1942 ();
 sky130_fd_sc_hd__decap_3 PHY_1943 ();
 sky130_fd_sc_hd__decap_3 PHY_1944 ();
 sky130_fd_sc_hd__decap_3 PHY_1945 ();
 sky130_fd_sc_hd__decap_3 PHY_1946 ();
 sky130_fd_sc_hd__decap_3 PHY_1947 ();
 sky130_fd_sc_hd__decap_3 PHY_1948 ();
 sky130_fd_sc_hd__decap_3 PHY_1949 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_1950 ();
 sky130_fd_sc_hd__decap_3 PHY_1951 ();
 sky130_fd_sc_hd__decap_3 PHY_1952 ();
 sky130_fd_sc_hd__decap_3 PHY_1953 ();
 sky130_fd_sc_hd__decap_3 PHY_1954 ();
 sky130_fd_sc_hd__decap_3 PHY_1955 ();
 sky130_fd_sc_hd__decap_3 PHY_1956 ();
 sky130_fd_sc_hd__decap_3 PHY_1957 ();
 sky130_fd_sc_hd__decap_3 PHY_1958 ();
 sky130_fd_sc_hd__decap_3 PHY_1959 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_1960 ();
 sky130_fd_sc_hd__decap_3 PHY_1961 ();
 sky130_fd_sc_hd__decap_3 PHY_1962 ();
 sky130_fd_sc_hd__decap_3 PHY_1963 ();
 sky130_fd_sc_hd__decap_3 PHY_1964 ();
 sky130_fd_sc_hd__decap_3 PHY_1965 ();
 sky130_fd_sc_hd__decap_3 PHY_1966 ();
 sky130_fd_sc_hd__decap_3 PHY_1967 ();
 sky130_fd_sc_hd__decap_3 PHY_1968 ();
 sky130_fd_sc_hd__decap_3 PHY_1969 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_1970 ();
 sky130_fd_sc_hd__decap_3 PHY_1971 ();
 sky130_fd_sc_hd__decap_3 PHY_1972 ();
 sky130_fd_sc_hd__decap_3 PHY_1973 ();
 sky130_fd_sc_hd__decap_3 PHY_1974 ();
 sky130_fd_sc_hd__decap_3 PHY_1975 ();
 sky130_fd_sc_hd__decap_3 PHY_1976 ();
 sky130_fd_sc_hd__decap_3 PHY_1977 ();
 sky130_fd_sc_hd__decap_3 PHY_1978 ();
 sky130_fd_sc_hd__decap_3 PHY_1979 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_1980 ();
 sky130_fd_sc_hd__decap_3 PHY_1981 ();
 sky130_fd_sc_hd__decap_3 PHY_1982 ();
 sky130_fd_sc_hd__decap_3 PHY_1983 ();
 sky130_fd_sc_hd__decap_3 PHY_1984 ();
 sky130_fd_sc_hd__decap_3 PHY_1985 ();
 sky130_fd_sc_hd__decap_3 PHY_1986 ();
 sky130_fd_sc_hd__decap_3 PHY_1987 ();
 sky130_fd_sc_hd__decap_3 PHY_1988 ();
 sky130_fd_sc_hd__decap_3 PHY_1989 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_1990 ();
 sky130_fd_sc_hd__decap_3 PHY_1991 ();
 sky130_fd_sc_hd__decap_3 PHY_1992 ();
 sky130_fd_sc_hd__decap_3 PHY_1993 ();
 sky130_fd_sc_hd__decap_3 PHY_1994 ();
 sky130_fd_sc_hd__decap_3 PHY_1995 ();
 sky130_fd_sc_hd__decap_3 PHY_1996 ();
 sky130_fd_sc_hd__decap_3 PHY_1997 ();
 sky130_fd_sc_hd__decap_3 PHY_1998 ();
 sky130_fd_sc_hd__decap_3 PHY_1999 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_2000 ();
 sky130_fd_sc_hd__decap_3 PHY_2001 ();
 sky130_fd_sc_hd__decap_3 PHY_2002 ();
 sky130_fd_sc_hd__decap_3 PHY_2003 ();
 sky130_fd_sc_hd__decap_3 PHY_2004 ();
 sky130_fd_sc_hd__decap_3 PHY_2005 ();
 sky130_fd_sc_hd__decap_3 PHY_2006 ();
 sky130_fd_sc_hd__decap_3 PHY_2007 ();
 sky130_fd_sc_hd__decap_3 PHY_2008 ();
 sky130_fd_sc_hd__decap_3 PHY_2009 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_2010 ();
 sky130_fd_sc_hd__decap_3 PHY_2011 ();
 sky130_fd_sc_hd__decap_3 PHY_2012 ();
 sky130_fd_sc_hd__decap_3 PHY_2013 ();
 sky130_fd_sc_hd__decap_3 PHY_2014 ();
 sky130_fd_sc_hd__decap_3 PHY_2015 ();
 sky130_fd_sc_hd__decap_3 PHY_2016 ();
 sky130_fd_sc_hd__decap_3 PHY_2017 ();
 sky130_fd_sc_hd__decap_3 PHY_2018 ();
 sky130_fd_sc_hd__decap_3 PHY_2019 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_2020 ();
 sky130_fd_sc_hd__decap_3 PHY_2021 ();
 sky130_fd_sc_hd__decap_3 PHY_2022 ();
 sky130_fd_sc_hd__decap_3 PHY_2023 ();
 sky130_fd_sc_hd__decap_3 PHY_2024 ();
 sky130_fd_sc_hd__decap_3 PHY_2025 ();
 sky130_fd_sc_hd__decap_3 PHY_2026 ();
 sky130_fd_sc_hd__decap_3 PHY_2027 ();
 sky130_fd_sc_hd__decap_3 PHY_2028 ();
 sky130_fd_sc_hd__decap_3 PHY_2029 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_2030 ();
 sky130_fd_sc_hd__decap_3 PHY_2031 ();
 sky130_fd_sc_hd__decap_3 PHY_2032 ();
 sky130_fd_sc_hd__decap_3 PHY_2033 ();
 sky130_fd_sc_hd__decap_3 PHY_2034 ();
 sky130_fd_sc_hd__decap_3 PHY_2035 ();
 sky130_fd_sc_hd__decap_3 PHY_2036 ();
 sky130_fd_sc_hd__decap_3 PHY_2037 ();
 sky130_fd_sc_hd__decap_3 PHY_2038 ();
 sky130_fd_sc_hd__decap_3 PHY_2039 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_2040 ();
 sky130_fd_sc_hd__decap_3 PHY_2041 ();
 sky130_fd_sc_hd__decap_3 PHY_2042 ();
 sky130_fd_sc_hd__decap_3 PHY_2043 ();
 sky130_fd_sc_hd__decap_3 PHY_2044 ();
 sky130_fd_sc_hd__decap_3 PHY_2045 ();
 sky130_fd_sc_hd__decap_3 PHY_2046 ();
 sky130_fd_sc_hd__decap_3 PHY_2047 ();
 sky130_fd_sc_hd__decap_3 PHY_2048 ();
 sky130_fd_sc_hd__decap_3 PHY_2049 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_2050 ();
 sky130_fd_sc_hd__decap_3 PHY_2051 ();
 sky130_fd_sc_hd__decap_3 PHY_2052 ();
 sky130_fd_sc_hd__decap_3 PHY_2053 ();
 sky130_fd_sc_hd__decap_3 PHY_2054 ();
 sky130_fd_sc_hd__decap_3 PHY_2055 ();
 sky130_fd_sc_hd__decap_3 PHY_2056 ();
 sky130_fd_sc_hd__decap_3 PHY_2057 ();
 sky130_fd_sc_hd__decap_3 PHY_2058 ();
 sky130_fd_sc_hd__decap_3 PHY_2059 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_2060 ();
 sky130_fd_sc_hd__decap_3 PHY_2061 ();
 sky130_fd_sc_hd__decap_3 PHY_2062 ();
 sky130_fd_sc_hd__decap_3 PHY_2063 ();
 sky130_fd_sc_hd__decap_3 PHY_2064 ();
 sky130_fd_sc_hd__decap_3 PHY_2065 ();
 sky130_fd_sc_hd__decap_3 PHY_2066 ();
 sky130_fd_sc_hd__decap_3 PHY_2067 ();
 sky130_fd_sc_hd__decap_3 PHY_2068 ();
 sky130_fd_sc_hd__decap_3 PHY_2069 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_2070 ();
 sky130_fd_sc_hd__decap_3 PHY_2071 ();
 sky130_fd_sc_hd__decap_3 PHY_2072 ();
 sky130_fd_sc_hd__decap_3 PHY_2073 ();
 sky130_fd_sc_hd__decap_3 PHY_2074 ();
 sky130_fd_sc_hd__decap_3 PHY_2075 ();
 sky130_fd_sc_hd__decap_3 PHY_2076 ();
 sky130_fd_sc_hd__decap_3 PHY_2077 ();
 sky130_fd_sc_hd__decap_3 PHY_2078 ();
 sky130_fd_sc_hd__decap_3 PHY_2079 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_2080 ();
 sky130_fd_sc_hd__decap_3 PHY_2081 ();
 sky130_fd_sc_hd__decap_3 PHY_2082 ();
 sky130_fd_sc_hd__decap_3 PHY_2083 ();
 sky130_fd_sc_hd__decap_3 PHY_2084 ();
 sky130_fd_sc_hd__decap_3 PHY_2085 ();
 sky130_fd_sc_hd__decap_3 PHY_2086 ();
 sky130_fd_sc_hd__decap_3 PHY_2087 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__decap_3 PHY_644 ();
 sky130_fd_sc_hd__decap_3 PHY_645 ();
 sky130_fd_sc_hd__decap_3 PHY_646 ();
 sky130_fd_sc_hd__decap_3 PHY_647 ();
 sky130_fd_sc_hd__decap_3 PHY_648 ();
 sky130_fd_sc_hd__decap_3 PHY_649 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_650 ();
 sky130_fd_sc_hd__decap_3 PHY_651 ();
 sky130_fd_sc_hd__decap_3 PHY_652 ();
 sky130_fd_sc_hd__decap_3 PHY_653 ();
 sky130_fd_sc_hd__decap_3 PHY_654 ();
 sky130_fd_sc_hd__decap_3 PHY_655 ();
 sky130_fd_sc_hd__decap_3 PHY_656 ();
 sky130_fd_sc_hd__decap_3 PHY_657 ();
 sky130_fd_sc_hd__decap_3 PHY_658 ();
 sky130_fd_sc_hd__decap_3 PHY_659 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_660 ();
 sky130_fd_sc_hd__decap_3 PHY_661 ();
 sky130_fd_sc_hd__decap_3 PHY_662 ();
 sky130_fd_sc_hd__decap_3 PHY_663 ();
 sky130_fd_sc_hd__decap_3 PHY_664 ();
 sky130_fd_sc_hd__decap_3 PHY_665 ();
 sky130_fd_sc_hd__decap_3 PHY_666 ();
 sky130_fd_sc_hd__decap_3 PHY_667 ();
 sky130_fd_sc_hd__decap_3 PHY_668 ();
 sky130_fd_sc_hd__decap_3 PHY_669 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_670 ();
 sky130_fd_sc_hd__decap_3 PHY_671 ();
 sky130_fd_sc_hd__decap_3 PHY_672 ();
 sky130_fd_sc_hd__decap_3 PHY_673 ();
 sky130_fd_sc_hd__decap_3 PHY_674 ();
 sky130_fd_sc_hd__decap_3 PHY_675 ();
 sky130_fd_sc_hd__decap_3 PHY_676 ();
 sky130_fd_sc_hd__decap_3 PHY_677 ();
 sky130_fd_sc_hd__decap_3 PHY_678 ();
 sky130_fd_sc_hd__decap_3 PHY_679 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_680 ();
 sky130_fd_sc_hd__decap_3 PHY_681 ();
 sky130_fd_sc_hd__decap_3 PHY_682 ();
 sky130_fd_sc_hd__decap_3 PHY_683 ();
 sky130_fd_sc_hd__decap_3 PHY_684 ();
 sky130_fd_sc_hd__decap_3 PHY_685 ();
 sky130_fd_sc_hd__decap_3 PHY_686 ();
 sky130_fd_sc_hd__decap_3 PHY_687 ();
 sky130_fd_sc_hd__decap_3 PHY_688 ();
 sky130_fd_sc_hd__decap_3 PHY_689 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_690 ();
 sky130_fd_sc_hd__decap_3 PHY_691 ();
 sky130_fd_sc_hd__decap_3 PHY_692 ();
 sky130_fd_sc_hd__decap_3 PHY_693 ();
 sky130_fd_sc_hd__decap_3 PHY_694 ();
 sky130_fd_sc_hd__decap_3 PHY_695 ();
 sky130_fd_sc_hd__decap_3 PHY_696 ();
 sky130_fd_sc_hd__decap_3 PHY_697 ();
 sky130_fd_sc_hd__decap_3 PHY_698 ();
 sky130_fd_sc_hd__decap_3 PHY_699 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_700 ();
 sky130_fd_sc_hd__decap_3 PHY_701 ();
 sky130_fd_sc_hd__decap_3 PHY_702 ();
 sky130_fd_sc_hd__decap_3 PHY_703 ();
 sky130_fd_sc_hd__decap_3 PHY_704 ();
 sky130_fd_sc_hd__decap_3 PHY_705 ();
 sky130_fd_sc_hd__decap_3 PHY_706 ();
 sky130_fd_sc_hd__decap_3 PHY_707 ();
 sky130_fd_sc_hd__decap_3 PHY_708 ();
 sky130_fd_sc_hd__decap_3 PHY_709 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_710 ();
 sky130_fd_sc_hd__decap_3 PHY_711 ();
 sky130_fd_sc_hd__decap_3 PHY_712 ();
 sky130_fd_sc_hd__decap_3 PHY_713 ();
 sky130_fd_sc_hd__decap_3 PHY_714 ();
 sky130_fd_sc_hd__decap_3 PHY_715 ();
 sky130_fd_sc_hd__decap_3 PHY_716 ();
 sky130_fd_sc_hd__decap_3 PHY_717 ();
 sky130_fd_sc_hd__decap_3 PHY_718 ();
 sky130_fd_sc_hd__decap_3 PHY_719 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_720 ();
 sky130_fd_sc_hd__decap_3 PHY_721 ();
 sky130_fd_sc_hd__decap_3 PHY_722 ();
 sky130_fd_sc_hd__decap_3 PHY_723 ();
 sky130_fd_sc_hd__decap_3 PHY_724 ();
 sky130_fd_sc_hd__decap_3 PHY_725 ();
 sky130_fd_sc_hd__decap_3 PHY_726 ();
 sky130_fd_sc_hd__decap_3 PHY_727 ();
 sky130_fd_sc_hd__decap_3 PHY_728 ();
 sky130_fd_sc_hd__decap_3 PHY_729 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_730 ();
 sky130_fd_sc_hd__decap_3 PHY_731 ();
 sky130_fd_sc_hd__decap_3 PHY_732 ();
 sky130_fd_sc_hd__decap_3 PHY_733 ();
 sky130_fd_sc_hd__decap_3 PHY_734 ();
 sky130_fd_sc_hd__decap_3 PHY_735 ();
 sky130_fd_sc_hd__decap_3 PHY_736 ();
 sky130_fd_sc_hd__decap_3 PHY_737 ();
 sky130_fd_sc_hd__decap_3 PHY_738 ();
 sky130_fd_sc_hd__decap_3 PHY_739 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_740 ();
 sky130_fd_sc_hd__decap_3 PHY_741 ();
 sky130_fd_sc_hd__decap_3 PHY_742 ();
 sky130_fd_sc_hd__decap_3 PHY_743 ();
 sky130_fd_sc_hd__decap_3 PHY_744 ();
 sky130_fd_sc_hd__decap_3 PHY_745 ();
 sky130_fd_sc_hd__decap_3 PHY_746 ();
 sky130_fd_sc_hd__decap_3 PHY_747 ();
 sky130_fd_sc_hd__decap_3 PHY_748 ();
 sky130_fd_sc_hd__decap_3 PHY_749 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_750 ();
 sky130_fd_sc_hd__decap_3 PHY_751 ();
 sky130_fd_sc_hd__decap_3 PHY_752 ();
 sky130_fd_sc_hd__decap_3 PHY_753 ();
 sky130_fd_sc_hd__decap_3 PHY_754 ();
 sky130_fd_sc_hd__decap_3 PHY_755 ();
 sky130_fd_sc_hd__decap_3 PHY_756 ();
 sky130_fd_sc_hd__decap_3 PHY_757 ();
 sky130_fd_sc_hd__decap_3 PHY_758 ();
 sky130_fd_sc_hd__decap_3 PHY_759 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_760 ();
 sky130_fd_sc_hd__decap_3 PHY_761 ();
 sky130_fd_sc_hd__decap_3 PHY_762 ();
 sky130_fd_sc_hd__decap_3 PHY_763 ();
 sky130_fd_sc_hd__decap_3 PHY_764 ();
 sky130_fd_sc_hd__decap_3 PHY_765 ();
 sky130_fd_sc_hd__decap_3 PHY_766 ();
 sky130_fd_sc_hd__decap_3 PHY_767 ();
 sky130_fd_sc_hd__decap_3 PHY_768 ();
 sky130_fd_sc_hd__decap_3 PHY_769 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_770 ();
 sky130_fd_sc_hd__decap_3 PHY_771 ();
 sky130_fd_sc_hd__decap_3 PHY_772 ();
 sky130_fd_sc_hd__decap_3 PHY_773 ();
 sky130_fd_sc_hd__decap_3 PHY_774 ();
 sky130_fd_sc_hd__decap_3 PHY_775 ();
 sky130_fd_sc_hd__decap_3 PHY_776 ();
 sky130_fd_sc_hd__decap_3 PHY_777 ();
 sky130_fd_sc_hd__decap_3 PHY_778 ();
 sky130_fd_sc_hd__decap_3 PHY_779 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_780 ();
 sky130_fd_sc_hd__decap_3 PHY_781 ();
 sky130_fd_sc_hd__decap_3 PHY_782 ();
 sky130_fd_sc_hd__decap_3 PHY_783 ();
 sky130_fd_sc_hd__decap_3 PHY_784 ();
 sky130_fd_sc_hd__decap_3 PHY_785 ();
 sky130_fd_sc_hd__decap_3 PHY_786 ();
 sky130_fd_sc_hd__decap_3 PHY_787 ();
 sky130_fd_sc_hd__decap_3 PHY_788 ();
 sky130_fd_sc_hd__decap_3 PHY_789 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_790 ();
 sky130_fd_sc_hd__decap_3 PHY_791 ();
 sky130_fd_sc_hd__decap_3 PHY_792 ();
 sky130_fd_sc_hd__decap_3 PHY_793 ();
 sky130_fd_sc_hd__decap_3 PHY_794 ();
 sky130_fd_sc_hd__decap_3 PHY_795 ();
 sky130_fd_sc_hd__decap_3 PHY_796 ();
 sky130_fd_sc_hd__decap_3 PHY_797 ();
 sky130_fd_sc_hd__decap_3 PHY_798 ();
 sky130_fd_sc_hd__decap_3 PHY_799 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_800 ();
 sky130_fd_sc_hd__decap_3 PHY_801 ();
 sky130_fd_sc_hd__decap_3 PHY_802 ();
 sky130_fd_sc_hd__decap_3 PHY_803 ();
 sky130_fd_sc_hd__decap_3 PHY_804 ();
 sky130_fd_sc_hd__decap_3 PHY_805 ();
 sky130_fd_sc_hd__decap_3 PHY_806 ();
 sky130_fd_sc_hd__decap_3 PHY_807 ();
 sky130_fd_sc_hd__decap_3 PHY_808 ();
 sky130_fd_sc_hd__decap_3 PHY_809 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_810 ();
 sky130_fd_sc_hd__decap_3 PHY_811 ();
 sky130_fd_sc_hd__decap_3 PHY_812 ();
 sky130_fd_sc_hd__decap_3 PHY_813 ();
 sky130_fd_sc_hd__decap_3 PHY_814 ();
 sky130_fd_sc_hd__decap_3 PHY_815 ();
 sky130_fd_sc_hd__decap_3 PHY_816 ();
 sky130_fd_sc_hd__decap_3 PHY_817 ();
 sky130_fd_sc_hd__decap_3 PHY_818 ();
 sky130_fd_sc_hd__decap_3 PHY_819 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_820 ();
 sky130_fd_sc_hd__decap_3 PHY_821 ();
 sky130_fd_sc_hd__decap_3 PHY_822 ();
 sky130_fd_sc_hd__decap_3 PHY_823 ();
 sky130_fd_sc_hd__decap_3 PHY_824 ();
 sky130_fd_sc_hd__decap_3 PHY_825 ();
 sky130_fd_sc_hd__decap_3 PHY_826 ();
 sky130_fd_sc_hd__decap_3 PHY_827 ();
 sky130_fd_sc_hd__decap_3 PHY_828 ();
 sky130_fd_sc_hd__decap_3 PHY_829 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_830 ();
 sky130_fd_sc_hd__decap_3 PHY_831 ();
 sky130_fd_sc_hd__decap_3 PHY_832 ();
 sky130_fd_sc_hd__decap_3 PHY_833 ();
 sky130_fd_sc_hd__decap_3 PHY_834 ();
 sky130_fd_sc_hd__decap_3 PHY_835 ();
 sky130_fd_sc_hd__decap_3 PHY_836 ();
 sky130_fd_sc_hd__decap_3 PHY_837 ();
 sky130_fd_sc_hd__decap_3 PHY_838 ();
 sky130_fd_sc_hd__decap_3 PHY_839 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_840 ();
 sky130_fd_sc_hd__decap_3 PHY_841 ();
 sky130_fd_sc_hd__decap_3 PHY_842 ();
 sky130_fd_sc_hd__decap_3 PHY_843 ();
 sky130_fd_sc_hd__decap_3 PHY_844 ();
 sky130_fd_sc_hd__decap_3 PHY_845 ();
 sky130_fd_sc_hd__decap_3 PHY_846 ();
 sky130_fd_sc_hd__decap_3 PHY_847 ();
 sky130_fd_sc_hd__decap_3 PHY_848 ();
 sky130_fd_sc_hd__decap_3 PHY_849 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_850 ();
 sky130_fd_sc_hd__decap_3 PHY_851 ();
 sky130_fd_sc_hd__decap_3 PHY_852 ();
 sky130_fd_sc_hd__decap_3 PHY_853 ();
 sky130_fd_sc_hd__decap_3 PHY_854 ();
 sky130_fd_sc_hd__decap_3 PHY_855 ();
 sky130_fd_sc_hd__decap_3 PHY_856 ();
 sky130_fd_sc_hd__decap_3 PHY_857 ();
 sky130_fd_sc_hd__decap_3 PHY_858 ();
 sky130_fd_sc_hd__decap_3 PHY_859 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_860 ();
 sky130_fd_sc_hd__decap_3 PHY_861 ();
 sky130_fd_sc_hd__decap_3 PHY_862 ();
 sky130_fd_sc_hd__decap_3 PHY_863 ();
 sky130_fd_sc_hd__decap_3 PHY_864 ();
 sky130_fd_sc_hd__decap_3 PHY_865 ();
 sky130_fd_sc_hd__decap_3 PHY_866 ();
 sky130_fd_sc_hd__decap_3 PHY_867 ();
 sky130_fd_sc_hd__decap_3 PHY_868 ();
 sky130_fd_sc_hd__decap_3 PHY_869 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_870 ();
 sky130_fd_sc_hd__decap_3 PHY_871 ();
 sky130_fd_sc_hd__decap_3 PHY_872 ();
 sky130_fd_sc_hd__decap_3 PHY_873 ();
 sky130_fd_sc_hd__decap_3 PHY_874 ();
 sky130_fd_sc_hd__decap_3 PHY_875 ();
 sky130_fd_sc_hd__decap_3 PHY_876 ();
 sky130_fd_sc_hd__decap_3 PHY_877 ();
 sky130_fd_sc_hd__decap_3 PHY_878 ();
 sky130_fd_sc_hd__decap_3 PHY_879 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_880 ();
 sky130_fd_sc_hd__decap_3 PHY_881 ();
 sky130_fd_sc_hd__decap_3 PHY_882 ();
 sky130_fd_sc_hd__decap_3 PHY_883 ();
 sky130_fd_sc_hd__decap_3 PHY_884 ();
 sky130_fd_sc_hd__decap_3 PHY_885 ();
 sky130_fd_sc_hd__decap_3 PHY_886 ();
 sky130_fd_sc_hd__decap_3 PHY_887 ();
 sky130_fd_sc_hd__decap_3 PHY_888 ();
 sky130_fd_sc_hd__decap_3 PHY_889 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_890 ();
 sky130_fd_sc_hd__decap_3 PHY_891 ();
 sky130_fd_sc_hd__decap_3 PHY_892 ();
 sky130_fd_sc_hd__decap_3 PHY_893 ();
 sky130_fd_sc_hd__decap_3 PHY_894 ();
 sky130_fd_sc_hd__decap_3 PHY_895 ();
 sky130_fd_sc_hd__decap_3 PHY_896 ();
 sky130_fd_sc_hd__decap_3 PHY_897 ();
 sky130_fd_sc_hd__decap_3 PHY_898 ();
 sky130_fd_sc_hd__decap_3 PHY_899 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_900 ();
 sky130_fd_sc_hd__decap_3 PHY_901 ();
 sky130_fd_sc_hd__decap_3 PHY_902 ();
 sky130_fd_sc_hd__decap_3 PHY_903 ();
 sky130_fd_sc_hd__decap_3 PHY_904 ();
 sky130_fd_sc_hd__decap_3 PHY_905 ();
 sky130_fd_sc_hd__decap_3 PHY_906 ();
 sky130_fd_sc_hd__decap_3 PHY_907 ();
 sky130_fd_sc_hd__decap_3 PHY_908 ();
 sky130_fd_sc_hd__decap_3 PHY_909 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_910 ();
 sky130_fd_sc_hd__decap_3 PHY_911 ();
 sky130_fd_sc_hd__decap_3 PHY_912 ();
 sky130_fd_sc_hd__decap_3 PHY_913 ();
 sky130_fd_sc_hd__decap_3 PHY_914 ();
 sky130_fd_sc_hd__decap_3 PHY_915 ();
 sky130_fd_sc_hd__decap_3 PHY_916 ();
 sky130_fd_sc_hd__decap_3 PHY_917 ();
 sky130_fd_sc_hd__decap_3 PHY_918 ();
 sky130_fd_sc_hd__decap_3 PHY_919 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_920 ();
 sky130_fd_sc_hd__decap_3 PHY_921 ();
 sky130_fd_sc_hd__decap_3 PHY_922 ();
 sky130_fd_sc_hd__decap_3 PHY_923 ();
 sky130_fd_sc_hd__decap_3 PHY_924 ();
 sky130_fd_sc_hd__decap_3 PHY_925 ();
 sky130_fd_sc_hd__decap_3 PHY_926 ();
 sky130_fd_sc_hd__decap_3 PHY_927 ();
 sky130_fd_sc_hd__decap_3 PHY_928 ();
 sky130_fd_sc_hd__decap_3 PHY_929 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_930 ();
 sky130_fd_sc_hd__decap_3 PHY_931 ();
 sky130_fd_sc_hd__decap_3 PHY_932 ();
 sky130_fd_sc_hd__decap_3 PHY_933 ();
 sky130_fd_sc_hd__decap_3 PHY_934 ();
 sky130_fd_sc_hd__decap_3 PHY_935 ();
 sky130_fd_sc_hd__decap_3 PHY_936 ();
 sky130_fd_sc_hd__decap_3 PHY_937 ();
 sky130_fd_sc_hd__decap_3 PHY_938 ();
 sky130_fd_sc_hd__decap_3 PHY_939 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_940 ();
 sky130_fd_sc_hd__decap_3 PHY_941 ();
 sky130_fd_sc_hd__decap_3 PHY_942 ();
 sky130_fd_sc_hd__decap_3 PHY_943 ();
 sky130_fd_sc_hd__decap_3 PHY_944 ();
 sky130_fd_sc_hd__decap_3 PHY_945 ();
 sky130_fd_sc_hd__decap_3 PHY_946 ();
 sky130_fd_sc_hd__decap_3 PHY_947 ();
 sky130_fd_sc_hd__decap_3 PHY_948 ();
 sky130_fd_sc_hd__decap_3 PHY_949 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_950 ();
 sky130_fd_sc_hd__decap_3 PHY_951 ();
 sky130_fd_sc_hd__decap_3 PHY_952 ();
 sky130_fd_sc_hd__decap_3 PHY_953 ();
 sky130_fd_sc_hd__decap_3 PHY_954 ();
 sky130_fd_sc_hd__decap_3 PHY_955 ();
 sky130_fd_sc_hd__decap_3 PHY_956 ();
 sky130_fd_sc_hd__decap_3 PHY_957 ();
 sky130_fd_sc_hd__decap_3 PHY_958 ();
 sky130_fd_sc_hd__decap_3 PHY_959 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_960 ();
 sky130_fd_sc_hd__decap_3 PHY_961 ();
 sky130_fd_sc_hd__decap_3 PHY_962 ();
 sky130_fd_sc_hd__decap_3 PHY_963 ();
 sky130_fd_sc_hd__decap_3 PHY_964 ();
 sky130_fd_sc_hd__decap_3 PHY_965 ();
 sky130_fd_sc_hd__decap_3 PHY_966 ();
 sky130_fd_sc_hd__decap_3 PHY_967 ();
 sky130_fd_sc_hd__decap_3 PHY_968 ();
 sky130_fd_sc_hd__decap_3 PHY_969 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_970 ();
 sky130_fd_sc_hd__decap_3 PHY_971 ();
 sky130_fd_sc_hd__decap_3 PHY_972 ();
 sky130_fd_sc_hd__decap_3 PHY_973 ();
 sky130_fd_sc_hd__decap_3 PHY_974 ();
 sky130_fd_sc_hd__decap_3 PHY_975 ();
 sky130_fd_sc_hd__decap_3 PHY_976 ();
 sky130_fd_sc_hd__decap_3 PHY_977 ();
 sky130_fd_sc_hd__decap_3 PHY_978 ();
 sky130_fd_sc_hd__decap_3 PHY_979 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_980 ();
 sky130_fd_sc_hd__decap_3 PHY_981 ();
 sky130_fd_sc_hd__decap_3 PHY_982 ();
 sky130_fd_sc_hd__decap_3 PHY_983 ();
 sky130_fd_sc_hd__decap_3 PHY_984 ();
 sky130_fd_sc_hd__decap_3 PHY_985 ();
 sky130_fd_sc_hd__decap_3 PHY_986 ();
 sky130_fd_sc_hd__decap_3 PHY_987 ();
 sky130_fd_sc_hd__decap_3 PHY_988 ();
 sky130_fd_sc_hd__decap_3 PHY_989 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_990 ();
 sky130_fd_sc_hd__decap_3 PHY_991 ();
 sky130_fd_sc_hd__decap_3 PHY_992 ();
 sky130_fd_sc_hd__decap_3 PHY_993 ();
 sky130_fd_sc_hd__decap_3 PHY_994 ();
 sky130_fd_sc_hd__decap_3 PHY_995 ();
 sky130_fd_sc_hd__decap_3 PHY_996 ();
 sky130_fd_sc_hd__decap_3 PHY_997 ();
 sky130_fd_sc_hd__decap_3 PHY_998 ();
 sky130_fd_sc_hd__decap_3 PHY_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8822 ();
 core U_CORE (.clk(clknet_1_0__leaf_wb_clk_i),
    .o_mem_write_M(core_mem_write_M),
    .rst(net1),
    .i_instr_ID({net45,
    net51,
    net60,
    net64,
    net72,
    net75,
    net81,
    net87,
    net90,
    net95,
    net98,
    net102,
    net109,
    net112,
    net118,
    net124,
    net127,
    net131,
    net134,
    net138,
    net142,
    net147,
    net23,
    net25,
    net29,
    net32,
    net35,
    net38,
    net42,
    net57,
    net104,
    net150}),
    .i_read_data_M({net334,
    net363,
    net403,
    net338,
    \data_reg[27] ,
    \data_reg[26] ,
    \data_reg[25] ,
    \data_reg[24] ,
    \data_reg[23] ,
    net454,
    net463,
    \data_reg[20] ,
    net380,
    net460,
    net423,
    net418,
    \data_reg[15] ,
    net441,
    net433,
    net451,
    net401,
    net416,
    \data_reg[9] ,
    \data_reg[8] ,
    net161,
    net167,
    net170,
    net176,
    net182,
    net199,
    net259,
    net305}),
    .o_data_addr_M({\core_data_addr_M[31] ,
    \core_data_addr_M[30] ,
    \core_data_addr_M[29] ,
    \core_data_addr_M[28] ,
    \core_data_addr_M[27] ,
    \core_data_addr_M[26] ,
    \core_data_addr_M[25] ,
    \core_data_addr_M[24] ,
    \core_data_addr_M[23] ,
    \core_data_addr_M[22] ,
    \core_data_addr_M[21] ,
    \core_data_addr_M[20] ,
    \core_data_addr_M[19] ,
    \core_data_addr_M[18] ,
    \core_data_addr_M[17] ,
    \core_data_addr_M[16] ,
    \core_data_addr_M[15] ,
    \core_data_addr_M[14] ,
    \core_data_addr_M[13] ,
    \core_data_addr_M[12] ,
    \core_data_addr_M[11] ,
    \core_data_addr_M[10] ,
    \core_data_addr_M[9] ,
    \core_data_addr_M[8] ,
    \core_data_addr_M[7] ,
    \core_data_addr_M[6] ,
    \core_data_addr_M[5] ,
    \core_data_addr_M[4] ,
    \core_data_addr_M[3] ,
    \core_data_addr_M[2] ,
    \core_data_addr_M[1] ,
    \core_data_addr_M[0] }),
    .o_funct3_MEM({\funct3[2] ,
    \funct3[1] ,
    \funct3[0] }),
    .o_pc_IF({\core_pc_IF[31] ,
    \core_pc_IF[30] ,
    \core_pc_IF[29] ,
    \core_pc_IF[28] ,
    \core_pc_IF[27] ,
    \core_pc_IF[26] ,
    \core_pc_IF[25] ,
    \core_pc_IF[24] ,
    \core_pc_IF[23] ,
    \core_pc_IF[22] ,
    \core_pc_IF[21] ,
    \core_pc_IF[20] ,
    \core_pc_IF[19] ,
    \core_pc_IF[18] ,
    \core_pc_IF[17] ,
    \core_pc_IF[16] ,
    \core_pc_IF[15] ,
    \core_pc_IF[14] ,
    \core_pc_IF[13] ,
    \core_pc_IF[12] ,
    \core_pc_IF[11] ,
    \core_pc_IF[10] ,
    \core_pc_IF[9] ,
    \core_pc_IF[8] ,
    \core_pc_IF[7] ,
    \core_pc_IF[6] ,
    \core_pc_IF[5] ,
    \core_pc_IF[4] ,
    \core_pc_IF[3] ,
    \core_pc_IF[2] ,
    \core_pc_IF[1] ,
    \core_pc_IF[0] }),
    .o_write_data_M({\core_write_data_M[31] ,
    \core_write_data_M[30] ,
    \core_write_data_M[29] ,
    \core_write_data_M[28] ,
    \core_write_data_M[27] ,
    \core_write_data_M[26] ,
    \core_write_data_M[25] ,
    \core_write_data_M[24] ,
    \core_write_data_M[23] ,
    \core_write_data_M[22] ,
    \core_write_data_M[21] ,
    \core_write_data_M[20] ,
    \core_write_data_M[19] ,
    \core_write_data_M[18] ,
    \core_write_data_M[17] ,
    \core_write_data_M[16] ,
    \core_write_data_M[15] ,
    \core_write_data_M[14] ,
    \core_write_data_M[13] ,
    \core_write_data_M[12] ,
    \core_write_data_M[11] ,
    \core_write_data_M[10] ,
    \core_write_data_M[9] ,
    \core_write_data_M[8] ,
    \core_write_data_M[7] ,
    \core_write_data_M[6] ,
    \core_write_data_M[5] ,
    \core_write_data_M[4] ,
    \core_write_data_M[3] ,
    \core_write_data_M[2] ,
    \core_write_data_M[1] ,
    \core_write_data_M[0] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 U_DATA_MEM (.csb0(net313),
    .csb1(net323),
    .web0(write_sram_data_mem),
    .clk0(clknet_1_1__leaf_wb_clk_i),
    .clk1(net312),
    .addr0({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9}),
    .addr1({_NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16,
    _NC17,
    _NC18}),
    .din0({\shifted_data[31] ,
    \shifted_data[30] ,
    \shifted_data[29] ,
    \shifted_data[28] ,
    \shifted_data[27] ,
    \shifted_data[26] ,
    \shifted_data[25] ,
    \shifted_data[24] ,
    \shifted_data[23] ,
    \shifted_data[22] ,
    \shifted_data[21] ,
    \shifted_data[20] ,
    \shifted_data[19] ,
    \shifted_data[18] ,
    \shifted_data[17] ,
    \shifted_data[16] ,
    \shifted_data[15] ,
    \shifted_data[14] ,
    \shifted_data[13] ,
    \shifted_data[12] ,
    \shifted_data[11] ,
    \shifted_data[10] ,
    \shifted_data[9] ,
    \shifted_data[8] ,
    \shifted_data[7] ,
    \shifted_data[6] ,
    \shifted_data[5] ,
    \shifted_data[4] ,
    \shifted_data[3] ,
    \shifted_data[2] ,
    \shifted_data[1] ,
    \shifted_data[0] }),
    .dout0({\core_read_data_M[31] ,
    \core_read_data_M[30] ,
    \core_read_data_M[29] ,
    \core_read_data_M[28] ,
    \core_read_data_M[27] ,
    \core_read_data_M[26] ,
    \core_read_data_M[25] ,
    \core_read_data_M[24] ,
    \core_read_data_M[23] ,
    \core_read_data_M[22] ,
    \core_read_data_M[21] ,
    \core_read_data_M[20] ,
    \core_read_data_M[19] ,
    \core_read_data_M[18] ,
    \core_read_data_M[17] ,
    \core_read_data_M[16] ,
    \core_read_data_M[15] ,
    \core_read_data_M[14] ,
    \core_read_data_M[13] ,
    \core_read_data_M[12] ,
    \core_read_data_M[11] ,
    \core_read_data_M[10] ,
    \core_read_data_M[9] ,
    \core_read_data_M[8] ,
    \core_read_data_M[7] ,
    \core_read_data_M[6] ,
    \core_read_data_M[5] ,
    \core_read_data_M[4] ,
    \core_read_data_M[3] ,
    \core_read_data_M[2] ,
    \core_read_data_M[1] ,
    \core_read_data_M[0] }),
    .dout1({\dummy_data2[31] ,
    \dummy_data2[30] ,
    \dummy_data2[29] ,
    \dummy_data2[28] ,
    \dummy_data2[27] ,
    \dummy_data2[26] ,
    \dummy_data2[25] ,
    \dummy_data2[24] ,
    \dummy_data2[23] ,
    \dummy_data2[22] ,
    \dummy_data2[21] ,
    \dummy_data2[20] ,
    \dummy_data2[19] ,
    \dummy_data2[18] ,
    \dummy_data2[17] ,
    \dummy_data2[16] ,
    \dummy_data2[15] ,
    \dummy_data2[14] ,
    \dummy_data2[13] ,
    \dummy_data2[12] ,
    \dummy_data2[11] ,
    \dummy_data2[10] ,
    \dummy_data2[9] ,
    \dummy_data2[8] ,
    \dummy_data2[7] ,
    \dummy_data2[6] ,
    \dummy_data2[5] ,
    \dummy_data2[4] ,
    \dummy_data2[3] ,
    \dummy_data2[2] ,
    \dummy_data2[1] ,
    \dummy_data2[0] }),
    .wmask0({net374,
    net369,
    net381,
    net383}));
 sky130_fd_sc_hd__conb_1 U_DATA_MEM_312 (.LO(net312));
 sky130_fd_sc_hd__conb_1 U_DATA_MEM_313 (.LO(net313));
 sky130_fd_sc_hd__conb_1 U_DATA_MEM_323 (.HI(net323));
 sky130_sram_2kbyte_1rw1r_32x512_8 U_INST_MEM (.csb0(net315),
    .csb1(net324),
    .web0(write_sram_inst_mem),
    .clk0(clknet_1_0__leaf_wb_clk_i),
    .clk1(net314),
    .addr0({_NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26,
    _NC27}),
    .addr1({_NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32,
    _NC33,
    _NC34,
    _NC35,
    _NC36}),
    .din0({\inst_mem_dat_i[31] ,
    \inst_mem_dat_i[30] ,
    \inst_mem_dat_i[29] ,
    \inst_mem_dat_i[28] ,
    \inst_mem_dat_i[27] ,
    \inst_mem_dat_i[26] ,
    \inst_mem_dat_i[25] ,
    \inst_mem_dat_i[24] ,
    \inst_mem_dat_i[23] ,
    \inst_mem_dat_i[22] ,
    \inst_mem_dat_i[21] ,
    \inst_mem_dat_i[20] ,
    \inst_mem_dat_i[19] ,
    \inst_mem_dat_i[18] ,
    \inst_mem_dat_i[17] ,
    \inst_mem_dat_i[16] ,
    \inst_mem_dat_i[15] ,
    \inst_mem_dat_i[14] ,
    \inst_mem_dat_i[13] ,
    \inst_mem_dat_i[12] ,
    \inst_mem_dat_i[11] ,
    \inst_mem_dat_i[10] ,
    \inst_mem_dat_i[9] ,
    \inst_mem_dat_i[8] ,
    \inst_mem_dat_i[7] ,
    \inst_mem_dat_i[6] ,
    \inst_mem_dat_i[5] ,
    \inst_mem_dat_i[4] ,
    \inst_mem_dat_i[3] ,
    \inst_mem_dat_i[2] ,
    \inst_mem_dat_i[1] ,
    \inst_mem_dat_i[0] }),
    .dout0({\core_instr_ID[31] ,
    \core_instr_ID[30] ,
    \core_instr_ID[29] ,
    \core_instr_ID[28] ,
    \core_instr_ID[27] ,
    \core_instr_ID[26] ,
    \core_instr_ID[25] ,
    \core_instr_ID[24] ,
    \core_instr_ID[23] ,
    \core_instr_ID[22] ,
    \core_instr_ID[21] ,
    \core_instr_ID[20] ,
    \core_instr_ID[19] ,
    \core_instr_ID[18] ,
    \core_instr_ID[17] ,
    \core_instr_ID[16] ,
    \core_instr_ID[15] ,
    \core_instr_ID[14] ,
    \core_instr_ID[13] ,
    \core_instr_ID[12] ,
    \core_instr_ID[11] ,
    \core_instr_ID[10] ,
    \core_instr_ID[9] ,
    \core_instr_ID[8] ,
    \core_instr_ID[7] ,
    \core_instr_ID[6] ,
    \core_instr_ID[5] ,
    \core_instr_ID[4] ,
    \core_instr_ID[3] ,
    \core_instr_ID[2] ,
    \core_instr_ID[1] ,
    \core_instr_ID[0] }),
    .dout1({\dummy_data[31] ,
    \dummy_data[30] ,
    \dummy_data[29] ,
    \dummy_data[28] ,
    \dummy_data[27] ,
    \dummy_data[26] ,
    \dummy_data[25] ,
    \dummy_data[24] ,
    \dummy_data[23] ,
    \dummy_data[22] ,
    \dummy_data[21] ,
    \dummy_data[20] ,
    \dummy_data[19] ,
    \dummy_data[18] ,
    \dummy_data[17] ,
    \dummy_data[16] ,
    \dummy_data[15] ,
    \dummy_data[14] ,
    \dummy_data[13] ,
    \dummy_data[12] ,
    \dummy_data[11] ,
    \dummy_data[10] ,
    \dummy_data[9] ,
    \dummy_data[8] ,
    \dummy_data[7] ,
    \dummy_data[6] ,
    \dummy_data[5] ,
    \dummy_data[4] ,
    \dummy_data[3] ,
    \dummy_data[2] ,
    \dummy_data[1] ,
    \dummy_data[0] }),
    .wmask0({net328,
    net327,
    net326,
    net325}));
 sky130_fd_sc_hd__conb_1 U_INST_MEM_314 (.LO(net314));
 sky130_fd_sc_hd__conb_1 U_INST_MEM_315 (.LO(net315));
 sky130_fd_sc_hd__conb_1 U_INST_MEM_324 (.HI(net324));
 sky130_fd_sc_hd__conb_1 U_INST_MEM_325 (.HI(net325));
 sky130_fd_sc_hd__conb_1 U_INST_MEM_326 (.HI(net326));
 sky130_fd_sc_hd__conb_1 U_INST_MEM_327 (.HI(net327));
 sky130_fd_sc_hd__conb_1 U_INST_MEM_328 (.HI(net328));
 uart_wbs_bridge U_UART_WB_BRIDGE (.clk(clknet_1_0__leaf_wb_clk_i),
    .i_start_rx(net5),
    .i_uart_rx(net3),
    .o_uart_tx(o_uart_tx),
    .rst(net2),
    .wb_ack_i(net329),
    .wb_cyc_o(uart_wb_cyc_o),
    .wb_stb_o(uart_wb_stb_o),
    .wb_we_o(uart_wb_we_o),
    .wb_adr_o({_NC37,
    _NC38,
    _NC39,
    _NC40,
    _NC41,
    _NC42,
    _NC43,
    _NC44,
    _NC45,
    _NC46,
    _NC47,
    _NC48,
    _NC49,
    _NC50,
    _NC51,
    _NC52}),
    .wb_dat_i({\uart_wb_dat_i[31] ,
    \uart_wb_dat_i[30] ,
    \uart_wb_dat_i[29] ,
    \uart_wb_dat_i[28] ,
    \uart_wb_dat_i[27] ,
    \uart_wb_dat_i[26] ,
    \uart_wb_dat_i[25] ,
    \uart_wb_dat_i[24] ,
    \uart_wb_dat_i[23] ,
    \uart_wb_dat_i[22] ,
    \uart_wb_dat_i[21] ,
    \uart_wb_dat_i[20] ,
    \uart_wb_dat_i[19] ,
    \uart_wb_dat_i[18] ,
    \uart_wb_dat_i[17] ,
    \uart_wb_dat_i[16] ,
    \uart_wb_dat_i[15] ,
    \uart_wb_dat_i[14] ,
    \uart_wb_dat_i[13] ,
    \uart_wb_dat_i[12] ,
    \uart_wb_dat_i[11] ,
    \uart_wb_dat_i[10] ,
    \uart_wb_dat_i[9] ,
    \uart_wb_dat_i[8] ,
    \uart_wb_dat_i[7] ,
    \uart_wb_dat_i[6] ,
    \uart_wb_dat_i[5] ,
    \uart_wb_dat_i[4] ,
    \uart_wb_dat_i[3] ,
    \uart_wb_dat_i[2] ,
    \uart_wb_dat_i[1] ,
    \uart_wb_dat_i[0] }),
    .wb_dat_o({\inst_mem_dat_i[31] ,
    \inst_mem_dat_i[30] ,
    \inst_mem_dat_i[29] ,
    \inst_mem_dat_i[28] ,
    \inst_mem_dat_i[27] ,
    \inst_mem_dat_i[26] ,
    \inst_mem_dat_i[25] ,
    \inst_mem_dat_i[24] ,
    \inst_mem_dat_i[23] ,
    \inst_mem_dat_i[22] ,
    \inst_mem_dat_i[21] ,
    \inst_mem_dat_i[20] ,
    \inst_mem_dat_i[19] ,
    \inst_mem_dat_i[18] ,
    \inst_mem_dat_i[17] ,
    \inst_mem_dat_i[16] ,
    \inst_mem_dat_i[15] ,
    \inst_mem_dat_i[14] ,
    \inst_mem_dat_i[13] ,
    \inst_mem_dat_i[12] ,
    \inst_mem_dat_i[11] ,
    \inst_mem_dat_i[10] ,
    \inst_mem_dat_i[9] ,
    \inst_mem_dat_i[8] ,
    \inst_mem_dat_i[7] ,
    \inst_mem_dat_i[6] ,
    \inst_mem_dat_i[5] ,
    \inst_mem_dat_i[4] ,
    \inst_mem_dat_i[3] ,
    \inst_mem_dat_i[2] ,
    \inst_mem_dat_i[1] ,
    \inst_mem_dat_i[0] }));
 sky130_fd_sc_hd__conb_1 U_UART_WB_BRIDGE_329 (.HI(net329));
 sky130_fd_sc_hd__inv_2 _105_ (.A(uart_wb_we_o),
    .Y(_000_));
 sky130_fd_sc_hd__nor2_1 _106_ (.A(net373),
    .B(net382),
    .Y(_001_));
 sky130_fd_sc_hd__or2_1 _107_ (.A(net373),
    .B(net382),
    .X(_002_));
 sky130_fd_sc_hd__or2_1 _108_ (.A(net382),
    .B(net348),
    .X(_003_));
 sky130_fd_sc_hd__nor3b_1 _109_ (.A(net349),
    .B(net373),
    .C_N(net163),
    .Y(_004_));
 sky130_fd_sc_hd__a31o_1 _110_ (.A1(net348),
    .A2(net280),
    .A3(net361),
    .B1(net344),
    .X(_005_));
 sky130_fd_sc_hd__a21o_2 _111_ (.A1(net382),
    .A2(net208),
    .B1(net399),
    .X(\data_reg[28] ));
 sky130_fd_sc_hd__a21o_4 _112_ (.A1(net382),
    .A2(net204),
    .B1(net399),
    .X(\data_reg[29] ));
 sky130_fd_sc_hd__a21o_1 _113_ (.A1(net382),
    .A2(net194),
    .B1(net399),
    .X(\data_reg[30] ));
 sky130_fd_sc_hd__a32o_2 _114_ (.A1(net348),
    .A2(net280),
    .A3(net361),
    .B1(net187),
    .B2(net382),
    .X(\data_reg[31] ));
 sky130_fd_sc_hd__nand2b_4 _115_ (.A_N(net310),
    .B(uart_wb_stb_o),
    .Y(_006_));
 sky130_fd_sc_hd__mux2_1 _116_ (.A0(\uart_wb_adr_o[0] ),
    .A1(\core_pc_IF[0] ),
    .S(_006_),
    .X(\inst_mem_adr_i[0] ));
 sky130_fd_sc_hd__mux2_1 _117_ (.A0(\uart_wb_adr_o[1] ),
    .A1(\core_pc_IF[1] ),
    .S(_006_),
    .X(\inst_mem_adr_i[1] ));
 sky130_fd_sc_hd__mux2_1 _118_ (.A0(\uart_wb_adr_o[2] ),
    .A1(\core_pc_IF[2] ),
    .S(_006_),
    .X(\inst_mem_adr_i[2] ));
 sky130_fd_sc_hd__mux2_1 _119_ (.A0(\uart_wb_adr_o[3] ),
    .A1(\core_pc_IF[3] ),
    .S(_006_),
    .X(\inst_mem_adr_i[3] ));
 sky130_fd_sc_hd__mux2_1 _120_ (.A0(\uart_wb_adr_o[4] ),
    .A1(\core_pc_IF[4] ),
    .S(_006_),
    .X(\inst_mem_adr_i[4] ));
 sky130_fd_sc_hd__mux2_1 _121_ (.A0(\uart_wb_adr_o[5] ),
    .A1(\core_pc_IF[5] ),
    .S(_006_),
    .X(\inst_mem_adr_i[5] ));
 sky130_fd_sc_hd__mux2_1 _122_ (.A0(\uart_wb_adr_o[6] ),
    .A1(\core_pc_IF[6] ),
    .S(_006_),
    .X(\inst_mem_adr_i[6] ));
 sky130_fd_sc_hd__mux2_1 _123_ (.A0(\uart_wb_adr_o[7] ),
    .A1(\core_pc_IF[7] ),
    .S(_006_),
    .X(\inst_mem_adr_i[7] ));
 sky130_fd_sc_hd__nand2_8 _124_ (.A(net310),
    .B(uart_wb_stb_o),
    .Y(_007_));
 sky130_fd_sc_hd__mux2_1 _125_ (.A0(\uart_wb_adr_o[2] ),
    .A1(\core_data_addr_M[2] ),
    .S(_007_),
    .X(\data_mem_adr_i[2] ));
 sky130_fd_sc_hd__mux2_1 _126_ (.A0(\uart_wb_adr_o[3] ),
    .A1(\core_data_addr_M[3] ),
    .S(net21),
    .X(\data_mem_adr_i[3] ));
 sky130_fd_sc_hd__mux2_1 _127_ (.A0(\uart_wb_adr_o[4] ),
    .A1(\core_data_addr_M[4] ),
    .S(net20),
    .X(\data_mem_adr_i[4] ));
 sky130_fd_sc_hd__mux2_1 _128_ (.A0(\uart_wb_adr_o[5] ),
    .A1(\core_data_addr_M[5] ),
    .S(net21),
    .X(\data_mem_adr_i[5] ));
 sky130_fd_sc_hd__mux2_1 _129_ (.A0(\uart_wb_adr_o[6] ),
    .A1(\core_data_addr_M[6] ),
    .S(_007_),
    .X(\data_mem_adr_i[6] ));
 sky130_fd_sc_hd__mux2_1 _130_ (.A0(\uart_wb_adr_o[7] ),
    .A1(\core_data_addr_M[7] ),
    .S(_007_),
    .X(\data_mem_adr_i[7] ));
 sky130_fd_sc_hd__and3_1 _131_ (.A(net311),
    .B(uart_wb_stb_o),
    .C(\uart_wb_adr_o[1] ),
    .X(_008_));
 sky130_fd_sc_hd__a21oi_4 _132_ (.A1(\core_data_addr_M[1] ),
    .A2(net21),
    .B1(_008_),
    .Y(_009_));
 sky130_fd_sc_hd__and3_2 _133_ (.A(net311),
    .B(uart_wb_stb_o),
    .C(\uart_wb_adr_o[0] ),
    .X(_010_));
 sky130_fd_sc_hd__a21oi_4 _134_ (.A1(\core_data_addr_M[0] ),
    .A2(net21),
    .B1(_010_),
    .Y(_011_));
 sky130_fd_sc_hd__a221o_4 _135_ (.A1(net311),
    .A2(uart_wb_cyc_o),
    .B1(\funct3[0] ),
    .B2(\funct3[1] ),
    .C1(\funct3[2] ),
    .X(_012_));
 sky130_fd_sc_hd__a21o_4 _136_ (.A1(net15),
    .A2(net14),
    .B1(_012_),
    .X(\mux_funct3[0] ));
 sky130_fd_sc_hd__or3b_4 _137_ (.A(\funct3[1] ),
    .B(\funct3[2] ),
    .C_N(\funct3[0] ),
    .X(_013_));
 sky130_fd_sc_hd__or3b_4 _138_ (.A(\funct3[0] ),
    .B(\funct3[2] ),
    .C_N(\funct3[1] ),
    .X(_014_));
 sky130_fd_sc_hd__nand3_2 _139_ (.A(net12),
    .B(_013_),
    .C(_014_),
    .Y(_015_));
 sky130_fd_sc_hd__a21o_4 _140_ (.A1(net15),
    .A2(_015_),
    .B1(_012_),
    .X(\mux_funct3[1] ));
 sky130_fd_sc_hd__o21ai_2 _141_ (.A1(net12),
    .A2(_013_),
    .B1(_014_),
    .Y(_016_));
 sky130_fd_sc_hd__and2b_4 _142_ (.A_N(net16),
    .B(net14),
    .X(_017_));
 sky130_fd_sc_hd__a211o_4 _143_ (.A1(net16),
    .A2(_016_),
    .B1(_017_),
    .C1(_012_),
    .X(\mux_funct3[2] ));
 sky130_fd_sc_hd__a21oi_1 _144_ (.A1(net12),
    .A2(_013_),
    .B1(net17),
    .Y(_018_));
 sky130_fd_sc_hd__a2111o_4 _145_ (.A1(net311),
    .A2(uart_wb_cyc_o),
    .B1(\funct3[1] ),
    .C1(\funct3[2] ),
    .D1(_018_),
    .X(\mux_funct3[3] ));
 sky130_fd_sc_hd__mux2_4 _146_ (.A0(net152),
    .A1(net305),
    .S(net310),
    .X(\uart_wb_dat_i[0] ));
 sky130_fd_sc_hd__mux2_4 _147_ (.A0(net107),
    .A1(net256),
    .S(net309),
    .X(\uart_wb_dat_i[1] ));
 sky130_fd_sc_hd__mux2_2 _148_ (.A0(net58),
    .A1(net199),
    .S(net309),
    .X(\uart_wb_dat_i[2] ));
 sky130_fd_sc_hd__mux2_2 _149_ (.A0(net43),
    .A1(net183),
    .S(net310),
    .X(\uart_wb_dat_i[3] ));
 sky130_fd_sc_hd__mux2_2 _150_ (.A0(net41),
    .A1(net178),
    .S(net310),
    .X(\uart_wb_dat_i[4] ));
 sky130_fd_sc_hd__mux2_4 _151_ (.A0(net37),
    .A1(net172),
    .S(net311),
    .X(\uart_wb_dat_i[5] ));
 sky130_fd_sc_hd__mux2_8 _152_ (.A0(net34),
    .A1(net166),
    .S(net310),
    .X(\uart_wb_dat_i[6] ));
 sky130_fd_sc_hd__mux2_1 _153_ (.A0(net30),
    .A1(net161),
    .S(net309),
    .X(\uart_wb_dat_i[7] ));
 sky130_fd_sc_hd__mux2_8 _154_ (.A0(net28),
    .A1(net157),
    .S(net311),
    .X(\uart_wb_dat_i[8] ));
 sky130_fd_sc_hd__mux2_2 _155_ (.A0(net23),
    .A1(net153),
    .S(net309),
    .X(\uart_wb_dat_i[9] ));
 sky130_fd_sc_hd__mux2_4 _156_ (.A0(net148),
    .A1(net301),
    .S(net309),
    .X(\uart_wb_dat_i[10] ));
 sky130_fd_sc_hd__mux2_8 _157_ (.A0(net145),
    .A1(net297),
    .S(net311),
    .X(\uart_wb_dat_i[11] ));
 sky130_fd_sc_hd__mux2_4 _158_ (.A0(net140),
    .A1(net293),
    .S(net311),
    .X(\uart_wb_dat_i[12] ));
 sky130_fd_sc_hd__mux2_4 _159_ (.A0(net136),
    .A1(net289),
    .S(net309),
    .X(\uart_wb_dat_i[13] ));
 sky130_fd_sc_hd__mux2_4 _160_ (.A0(net132),
    .A1(net285),
    .S(net310),
    .X(\uart_wb_dat_i[14] ));
 sky130_fd_sc_hd__mux2_1 _161_ (.A0(net128),
    .A1(net279),
    .S(net309),
    .X(\uart_wb_dat_i[15] ));
 sky130_fd_sc_hd__mux2_4 _162_ (.A0(net125),
    .A1(net275),
    .S(net310),
    .X(\uart_wb_dat_i[16] ));
 sky130_fd_sc_hd__mux2_4 _163_ (.A0(net121),
    .A1(net270),
    .S(net311),
    .X(\uart_wb_dat_i[17] ));
 sky130_fd_sc_hd__mux2_4 _164_ (.A0(net115),
    .A1(net265),
    .S(net311),
    .X(\uart_wb_dat_i[18] ));
 sky130_fd_sc_hd__mux2_4 _165_ (.A0(net109),
    .A1(net260),
    .S(net309),
    .X(\uart_wb_dat_i[19] ));
 sky130_fd_sc_hd__mux2_4 _166_ (.A0(net102),
    .A1(net251),
    .S(net310),
    .X(\uart_wb_dat_i[20] ));
 sky130_fd_sc_hd__mux2_4 _167_ (.A0(net100),
    .A1(net246),
    .S(net309),
    .X(\uart_wb_dat_i[21] ));
 sky130_fd_sc_hd__mux2_1 _168_ (.A0(net95),
    .A1(net241),
    .S(net310),
    .X(\uart_wb_dat_i[22] ));
 sky130_fd_sc_hd__mux2_2 _169_ (.A0(net91),
    .A1(net235),
    .S(net310),
    .X(\uart_wb_dat_i[23] ));
 sky130_fd_sc_hd__mux2_8 _170_ (.A0(net87),
    .A1(net230),
    .S(net310),
    .X(\uart_wb_dat_i[24] ));
 sky130_fd_sc_hd__mux2_2 _171_ (.A0(net84),
    .A1(net224),
    .S(net309),
    .X(\uart_wb_dat_i[25] ));
 sky130_fd_sc_hd__mux2_2 _172_ (.A0(net78),
    .A1(net219),
    .S(net309),
    .X(\uart_wb_dat_i[26] ));
 sky130_fd_sc_hd__mux2_4 _173_ (.A0(net72),
    .A1(net214),
    .S(net309),
    .X(\uart_wb_dat_i[27] ));
 sky130_fd_sc_hd__mux2_4 _174_ (.A0(net68),
    .A1(net208),
    .S(net309),
    .X(\uart_wb_dat_i[28] ));
 sky130_fd_sc_hd__mux2_4 _175_ (.A0(net61),
    .A1(net203),
    .S(net309),
    .X(\uart_wb_dat_i[29] ));
 sky130_fd_sc_hd__mux2_2 _176_ (.A0(net53),
    .A1(net193),
    .S(net309),
    .X(\uart_wb_dat_i[30] ));
 sky130_fd_sc_hd__mux2_2 _177_ (.A0(net48),
    .A1(net187),
    .S(net309),
    .X(\uart_wb_dat_i[31] ));
 sky130_fd_sc_hd__a21o_4 _178_ (.A1(net158),
    .A2(net349),
    .B1(net375),
    .X(\data_reg[8] ));
 sky130_fd_sc_hd__a21o_4 _179_ (.A1(net154),
    .A2(net349),
    .B1(net375),
    .X(\data_reg[9] ));
 sky130_fd_sc_hd__a21o_2 _180_ (.A1(net301),
    .A2(net349),
    .B1(net344),
    .X(\data_reg[10] ));
 sky130_fd_sc_hd__a21o_2 _181_ (.A1(net297),
    .A2(net349),
    .B1(net344),
    .X(\data_reg[11] ));
 sky130_fd_sc_hd__a21o_4 _182_ (.A1(net294),
    .A2(net349),
    .B1(net375),
    .X(\data_reg[12] ));
 sky130_fd_sc_hd__a21o_1 _183_ (.A1(net290),
    .A2(net349),
    .B1(net344),
    .X(\data_reg[13] ));
 sky130_fd_sc_hd__a21o_4 _184_ (.A1(net286),
    .A2(net349),
    .B1(net375),
    .X(\data_reg[14] ));
 sky130_fd_sc_hd__a31o_4 _185_ (.A1(net281),
    .A2(net387),
    .A3(net349),
    .B1(net399),
    .X(\data_reg[15] ));
 sky130_fd_sc_hd__a21o_1 _186_ (.A1(net382),
    .A2(net276),
    .B1(net399),
    .X(\data_reg[16] ));
 sky130_fd_sc_hd__a21o_1 _187_ (.A1(net382),
    .A2(net272),
    .B1(net399),
    .X(\data_reg[17] ));
 sky130_fd_sc_hd__a21o_2 _188_ (.A1(net382),
    .A2(net266),
    .B1(net399),
    .X(\data_reg[18] ));
 sky130_fd_sc_hd__a21o_2 _189_ (.A1(net382),
    .A2(net260),
    .B1(net399),
    .X(\data_reg[19] ));
 sky130_fd_sc_hd__a21o_4 _190_ (.A1(net382),
    .A2(net252),
    .B1(net399),
    .X(\data_reg[20] ));
 sky130_fd_sc_hd__a21o_1 _191_ (.A1(net382),
    .A2(net247),
    .B1(net399),
    .X(\data_reg[21] ));
 sky130_fd_sc_hd__a21o_4 _192_ (.A1(net382),
    .A2(net242),
    .B1(net399),
    .X(\data_reg[22] ));
 sky130_fd_sc_hd__a21o_4 _193_ (.A1(net382),
    .A2(net235),
    .B1(net399),
    .X(\data_reg[23] ));
 sky130_fd_sc_hd__a21o_4 _194_ (.A1(net386),
    .A2(net231),
    .B1(net399),
    .X(\data_reg[24] ));
 sky130_fd_sc_hd__a21o_4 _195_ (.A1(net382),
    .A2(net225),
    .B1(net399),
    .X(\data_reg[25] ));
 sky130_fd_sc_hd__a21o_4 _196_ (.A1(net386),
    .A2(net220),
    .B1(net399),
    .X(\data_reg[26] ));
 sky130_fd_sc_hd__a21o_4 _197_ (.A1(net386),
    .A2(net215),
    .B1(net399),
    .X(\data_reg[27] ));
 sky130_fd_sc_hd__or2_2 _198_ (.A(_000_),
    .B(_006_),
    .X(write_sram_inst_mem));
 sky130_fd_sc_hd__mux2_8 _199_ (.A0(uart_wb_we_o),
    .A1(core_mem_write_M),
    .S(net19),
    .X(_019_));
 sky130_fd_sc_hd__inv_6 _200_ (.A(_019_),
    .Y(write_sram_data_mem));
 sky130_fd_sc_hd__mux2_8 _201_ (.A0(\inst_mem_dat_i[0] ),
    .A1(\core_write_data_M[0] ),
    .S(net19),
    .X(_020_));
 sky130_fd_sc_hd__and3_4 _202_ (.A(net15),
    .B(net14),
    .C(_020_),
    .X(\shifted_data[0] ));
 sky130_fd_sc_hd__mux2_8 _203_ (.A0(\inst_mem_dat_i[1] ),
    .A1(\core_write_data_M[1] ),
    .S(net19),
    .X(_021_));
 sky130_fd_sc_hd__and3_4 _204_ (.A(net15),
    .B(net14),
    .C(_021_),
    .X(\shifted_data[1] ));
 sky130_fd_sc_hd__mux2_8 _205_ (.A0(\inst_mem_dat_i[2] ),
    .A1(\core_write_data_M[2] ),
    .S(net19),
    .X(_022_));
 sky130_fd_sc_hd__and3_4 _206_ (.A(net15),
    .B(net14),
    .C(_022_),
    .X(\shifted_data[2] ));
 sky130_fd_sc_hd__mux2_8 _207_ (.A0(\inst_mem_dat_i[3] ),
    .A1(\core_write_data_M[3] ),
    .S(net19),
    .X(_023_));
 sky130_fd_sc_hd__and3_4 _208_ (.A(net15),
    .B(net14),
    .C(_023_),
    .X(\shifted_data[3] ));
 sky130_fd_sc_hd__mux2_8 _209_ (.A0(\inst_mem_dat_i[4] ),
    .A1(\core_write_data_M[4] ),
    .S(net21),
    .X(_024_));
 sky130_fd_sc_hd__and3_4 _210_ (.A(net15),
    .B(net14),
    .C(_024_),
    .X(\shifted_data[4] ));
 sky130_fd_sc_hd__mux2_4 _211_ (.A0(\inst_mem_dat_i[5] ),
    .A1(\core_write_data_M[5] ),
    .S(net19),
    .X(_025_));
 sky130_fd_sc_hd__and3_4 _212_ (.A(net15),
    .B(net14),
    .C(_025_),
    .X(\shifted_data[5] ));
 sky130_fd_sc_hd__mux2_4 _213_ (.A0(\inst_mem_dat_i[6] ),
    .A1(\core_write_data_M[6] ),
    .S(net21),
    .X(_026_));
 sky130_fd_sc_hd__and3_4 _214_ (.A(net15),
    .B(net14),
    .C(_026_),
    .X(\shifted_data[6] ));
 sky130_fd_sc_hd__mux2_8 _215_ (.A0(\inst_mem_dat_i[7] ),
    .A1(\core_write_data_M[7] ),
    .S(net19),
    .X(_027_));
 sky130_fd_sc_hd__and3_4 _216_ (.A(net15),
    .B(net14),
    .C(_027_),
    .X(\shifted_data[7] ));
 sky130_fd_sc_hd__mux2_4 _217_ (.A0(\inst_mem_dat_i[8] ),
    .A1(\core_write_data_M[8] ),
    .S(net19),
    .X(_028_));
 sky130_fd_sc_hd__mux2_2 _218_ (.A0(_020_),
    .A1(_028_),
    .S(net12),
    .X(_029_));
 sky130_fd_sc_hd__and2_4 _219_ (.A(net15),
    .B(_029_),
    .X(\shifted_data[8] ));
 sky130_fd_sc_hd__mux2_2 _220_ (.A0(\inst_mem_dat_i[9] ),
    .A1(\core_write_data_M[9] ),
    .S(net19),
    .X(_030_));
 sky130_fd_sc_hd__mux2_2 _221_ (.A0(_021_),
    .A1(_030_),
    .S(net14),
    .X(_031_));
 sky130_fd_sc_hd__and2_4 _222_ (.A(net15),
    .B(_031_),
    .X(\shifted_data[9] ));
 sky130_fd_sc_hd__mux2_2 _223_ (.A0(\inst_mem_dat_i[10] ),
    .A1(\core_write_data_M[10] ),
    .S(net20),
    .X(_032_));
 sky130_fd_sc_hd__mux2_2 _224_ (.A0(_022_),
    .A1(_032_),
    .S(net12),
    .X(_033_));
 sky130_fd_sc_hd__and2_4 _225_ (.A(net15),
    .B(_033_),
    .X(\shifted_data[10] ));
 sky130_fd_sc_hd__mux2_4 _226_ (.A0(\inst_mem_dat_i[11] ),
    .A1(\core_write_data_M[11] ),
    .S(net19),
    .X(_034_));
 sky130_fd_sc_hd__mux2_2 _227_ (.A0(_023_),
    .A1(_034_),
    .S(net12),
    .X(_035_));
 sky130_fd_sc_hd__and2_4 _228_ (.A(net15),
    .B(_035_),
    .X(\shifted_data[11] ));
 sky130_fd_sc_hd__mux2_2 _229_ (.A0(\inst_mem_dat_i[12] ),
    .A1(\core_write_data_M[12] ),
    .S(net20),
    .X(_036_));
 sky130_fd_sc_hd__mux2_2 _230_ (.A0(_024_),
    .A1(_036_),
    .S(net12),
    .X(_037_));
 sky130_fd_sc_hd__and2_4 _231_ (.A(net15),
    .B(_037_),
    .X(\shifted_data[12] ));
 sky130_fd_sc_hd__mux2_4 _232_ (.A0(\inst_mem_dat_i[13] ),
    .A1(\core_write_data_M[13] ),
    .S(net20),
    .X(_038_));
 sky130_fd_sc_hd__mux2_2 _233_ (.A0(_025_),
    .A1(_038_),
    .S(net12),
    .X(_039_));
 sky130_fd_sc_hd__and2_4 _234_ (.A(net15),
    .B(_039_),
    .X(\shifted_data[13] ));
 sky130_fd_sc_hd__mux2_4 _235_ (.A0(\inst_mem_dat_i[14] ),
    .A1(\core_write_data_M[14] ),
    .S(net19),
    .X(_040_));
 sky130_fd_sc_hd__mux2_2 _236_ (.A0(_026_),
    .A1(_040_),
    .S(net12),
    .X(_041_));
 sky130_fd_sc_hd__and2_4 _237_ (.A(net16),
    .B(_041_),
    .X(\shifted_data[14] ));
 sky130_fd_sc_hd__mux2_4 _238_ (.A0(\inst_mem_dat_i[15] ),
    .A1(\core_write_data_M[15] ),
    .S(net19),
    .X(_042_));
 sky130_fd_sc_hd__mux2_2 _239_ (.A0(_027_),
    .A1(_042_),
    .S(net12),
    .X(_043_));
 sky130_fd_sc_hd__and2_4 _240_ (.A(net16),
    .B(_043_),
    .X(\shifted_data[15] ));
 sky130_fd_sc_hd__mux2_2 _241_ (.A0(\inst_mem_dat_i[16] ),
    .A1(\core_write_data_M[16] ),
    .S(net20),
    .X(_044_));
 sky130_fd_sc_hd__mux2_2 _242_ (.A0(_028_),
    .A1(_044_),
    .S(net12),
    .X(_045_));
 sky130_fd_sc_hd__a22o_4 _243_ (.A1(_017_),
    .A2(_020_),
    .B1(_045_),
    .B2(net16),
    .X(\shifted_data[16] ));
 sky130_fd_sc_hd__mux2_4 _244_ (.A0(\inst_mem_dat_i[17] ),
    .A1(\core_write_data_M[17] ),
    .S(net19),
    .X(_046_));
 sky130_fd_sc_hd__mux2_2 _245_ (.A0(_030_),
    .A1(_046_),
    .S(net12),
    .X(_047_));
 sky130_fd_sc_hd__a22o_4 _246_ (.A1(_017_),
    .A2(_021_),
    .B1(_047_),
    .B2(net16),
    .X(\shifted_data[17] ));
 sky130_fd_sc_hd__mux2_2 _247_ (.A0(\inst_mem_dat_i[18] ),
    .A1(\core_write_data_M[18] ),
    .S(net20),
    .X(_048_));
 sky130_fd_sc_hd__mux2_2 _248_ (.A0(_032_),
    .A1(_048_),
    .S(net12),
    .X(_049_));
 sky130_fd_sc_hd__a22o_4 _249_ (.A1(_017_),
    .A2(_022_),
    .B1(_049_),
    .B2(net16),
    .X(\shifted_data[18] ));
 sky130_fd_sc_hd__mux2_2 _250_ (.A0(\inst_mem_dat_i[19] ),
    .A1(\core_write_data_M[19] ),
    .S(net20),
    .X(_050_));
 sky130_fd_sc_hd__mux2_2 _251_ (.A0(_034_),
    .A1(_050_),
    .S(net12),
    .X(_051_));
 sky130_fd_sc_hd__a22o_4 _252_ (.A1(_017_),
    .A2(_023_),
    .B1(_051_),
    .B2(net16),
    .X(\shifted_data[19] ));
 sky130_fd_sc_hd__mux2_4 _253_ (.A0(\inst_mem_dat_i[20] ),
    .A1(\core_write_data_M[20] ),
    .S(net19),
    .X(_052_));
 sky130_fd_sc_hd__mux2_2 _254_ (.A0(_036_),
    .A1(_052_),
    .S(net12),
    .X(_053_));
 sky130_fd_sc_hd__a22o_4 _255_ (.A1(_017_),
    .A2(_024_),
    .B1(_053_),
    .B2(net16),
    .X(\shifted_data[20] ));
 sky130_fd_sc_hd__mux2_4 _256_ (.A0(\inst_mem_dat_i[21] ),
    .A1(\core_write_data_M[21] ),
    .S(net19),
    .X(_054_));
 sky130_fd_sc_hd__mux2_2 _257_ (.A0(_038_),
    .A1(_054_),
    .S(net12),
    .X(_055_));
 sky130_fd_sc_hd__a22o_4 _258_ (.A1(_017_),
    .A2(_025_),
    .B1(_055_),
    .B2(net17),
    .X(\shifted_data[21] ));
 sky130_fd_sc_hd__mux2_2 _259_ (.A0(\inst_mem_dat_i[22] ),
    .A1(\core_write_data_M[22] ),
    .S(net20),
    .X(_056_));
 sky130_fd_sc_hd__mux2_2 _260_ (.A0(_040_),
    .A1(_056_),
    .S(net13),
    .X(_057_));
 sky130_fd_sc_hd__a22o_4 _261_ (.A1(_017_),
    .A2(_026_),
    .B1(_057_),
    .B2(net16),
    .X(\shifted_data[22] ));
 sky130_fd_sc_hd__mux2_4 _262_ (.A0(\inst_mem_dat_i[23] ),
    .A1(\core_write_data_M[23] ),
    .S(net20),
    .X(_058_));
 sky130_fd_sc_hd__mux2_2 _263_ (.A0(_042_),
    .A1(_058_),
    .S(net13),
    .X(_059_));
 sky130_fd_sc_hd__a22o_4 _264_ (.A1(_017_),
    .A2(_027_),
    .B1(_059_),
    .B2(net17),
    .X(\shifted_data[23] ));
 sky130_fd_sc_hd__mux2_2 _265_ (.A0(\inst_mem_dat_i[24] ),
    .A1(\core_write_data_M[24] ),
    .S(net20),
    .X(_060_));
 sky130_fd_sc_hd__mux2_2 _266_ (.A0(_044_),
    .A1(_060_),
    .S(net13),
    .X(_061_));
 sky130_fd_sc_hd__mux2_8 _267_ (.A0(_029_),
    .A1(_061_),
    .S(net16),
    .X(\shifted_data[24] ));
 sky130_fd_sc_hd__mux2_2 _268_ (.A0(\inst_mem_dat_i[25] ),
    .A1(\core_write_data_M[25] ),
    .S(net20),
    .X(_062_));
 sky130_fd_sc_hd__mux2_2 _269_ (.A0(_046_),
    .A1(_062_),
    .S(net13),
    .X(_063_));
 sky130_fd_sc_hd__mux2_8 _270_ (.A0(_031_),
    .A1(_063_),
    .S(net16),
    .X(\shifted_data[25] ));
 sky130_fd_sc_hd__mux2_2 _271_ (.A0(\inst_mem_dat_i[26] ),
    .A1(\core_write_data_M[26] ),
    .S(net19),
    .X(_064_));
 sky130_fd_sc_hd__mux2_2 _272_ (.A0(_048_),
    .A1(_064_),
    .S(net13),
    .X(_065_));
 sky130_fd_sc_hd__mux2_8 _273_ (.A0(_033_),
    .A1(_065_),
    .S(net16),
    .X(\shifted_data[26] ));
 sky130_fd_sc_hd__mux2_2 _274_ (.A0(\inst_mem_dat_i[27] ),
    .A1(\core_write_data_M[27] ),
    .S(net20),
    .X(_066_));
 sky130_fd_sc_hd__mux2_2 _275_ (.A0(_050_),
    .A1(_066_),
    .S(net13),
    .X(_067_));
 sky130_fd_sc_hd__mux2_8 _276_ (.A0(_035_),
    .A1(_067_),
    .S(net16),
    .X(\shifted_data[27] ));
 sky130_fd_sc_hd__mux2_2 _277_ (.A0(\inst_mem_dat_i[28] ),
    .A1(\core_write_data_M[28] ),
    .S(net20),
    .X(_068_));
 sky130_fd_sc_hd__mux2_2 _278_ (.A0(_052_),
    .A1(_068_),
    .S(net13),
    .X(_069_));
 sky130_fd_sc_hd__mux2_8 _279_ (.A0(_037_),
    .A1(_069_),
    .S(net17),
    .X(\shifted_data[28] ));
 sky130_fd_sc_hd__mux2_2 _280_ (.A0(\inst_mem_dat_i[29] ),
    .A1(\core_write_data_M[29] ),
    .S(net20),
    .X(_070_));
 sky130_fd_sc_hd__mux2_4 _281_ (.A0(_054_),
    .A1(_070_),
    .S(net13),
    .X(_071_));
 sky130_fd_sc_hd__mux2_8 _282_ (.A0(_039_),
    .A1(_071_),
    .S(net17),
    .X(\shifted_data[29] ));
 sky130_fd_sc_hd__mux2_2 _283_ (.A0(\inst_mem_dat_i[30] ),
    .A1(\core_write_data_M[30] ),
    .S(net20),
    .X(_072_));
 sky130_fd_sc_hd__mux2_2 _284_ (.A0(_056_),
    .A1(_072_),
    .S(net13),
    .X(_073_));
 sky130_fd_sc_hd__mux2_8 _285_ (.A0(_041_),
    .A1(_073_),
    .S(net17),
    .X(\shifted_data[30] ));
 sky130_fd_sc_hd__mux2_2 _286_ (.A0(\inst_mem_dat_i[31] ),
    .A1(\core_write_data_M[31] ),
    .S(net21),
    .X(_074_));
 sky130_fd_sc_hd__mux2_4 _287_ (.A0(_058_),
    .A1(_074_),
    .S(net13),
    .X(_075_));
 sky130_fd_sc_hd__mux2_8 _288_ (.A0(_043_),
    .A1(_075_),
    .S(net17),
    .X(\shifted_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _289_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(\funct3[0] ),
    .Q(\funct3_s2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _290_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(\funct3[1] ),
    .Q(\funct3_s2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _291_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(\funct3[2] ),
    .Q(\funct3_s2[2] ));
 sky130_fd_sc_hd__clkbuf_2 _328_ (.A(o_uart_tx),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 _329_ (.A(o_uart_tx),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__buf_6 fanout12 (.A(net13),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_8 fanout13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_8 fanout14 (.A(_011_),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_8 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__buf_8 fanout16 (.A(net17),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_8 fanout17 (.A(_009_),
    .X(net17));
 sky130_fd_sc_hd__buf_12 fanout19 (.A(net20),
    .X(net19));
 sky130_fd_sc_hd__buf_8 fanout20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__buf_8 fanout21 (.A(_007_),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 fanout22 (.A(net386),
    .X(net22));
 sky130_fd_sc_hd__buf_8 fanout309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__buf_8 fanout310 (.A(net311),
    .X(net310));
 sky130_fd_sc_hd__buf_8 fanout311 (.A(net4),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net351),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net365),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\data_reg[11] ),
    .X(net438));
 sky130_fd_sc_hd__buf_1 hold104 (.A(net396),
    .X(net433));
 sky130_fd_sc_hd__buf_6 hold107 (.A(net479),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net347),
    .X(net340));
 sky130_fd_sc_hd__buf_4 hold117 (.A(\data_reg[12] ),
    .X(net451));
 sky130_fd_sc_hd__buf_6 hold12 (.A(_005_),
    .X(net341));
 sky130_fd_sc_hd__buf_6 hold120 (.A(\data_reg[22] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\data_reg[18] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\data_reg[21] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net371),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\data_reg[28] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net358),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\data_reg[14] ),
    .X(net479));
 sky130_fd_sc_hd__buf_2 hold15 (.A(net394),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net364),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net366),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net368),
    .X(net347));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold19 (.A(net340),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net367),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_8 hold20 (.A(_003_),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net385),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net335),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net330),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net336),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net22),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_2 hold26 (.A(net337),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net391),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net372),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net332),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net357),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net343),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_001_),
    .X(net360));
 sky130_fd_sc_hd__buf_1 hold32 (.A(net333),
    .X(net361));
 sky130_fd_sc_hd__buf_8 hold33 (.A(net341),
    .X(net362));
 sky130_fd_sc_hd__buf_8 hold34 (.A(\data_reg[30] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net397),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net345),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net339),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net346),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net331),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net360),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\funct3_s2[1] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net390),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net356),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net342),
    .X(net372));
 sky130_fd_sc_hd__buf_1 hold44 (.A(net359),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net378),
    .X(net386));
 sky130_fd_sc_hd__buf_2 hold46 (.A(net18),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net353),
    .X(net376));
 sky130_fd_sc_hd__buf_6 hold48 (.A(net355),
    .X(net377));
 sky130_fd_sc_hd__buf_2 hold49 (.A(net376),
    .X(net378));
 sky130_fd_sc_hd__buf_2 hold5 (.A(net419),
    .X(net334));
 sky130_fd_sc_hd__buf_6 hold50 (.A(net377),
    .X(net379));
 sky130_fd_sc_hd__buf_4 hold51 (.A(\data_reg[19] ),
    .X(net380));
 sky130_fd_sc_hd__buf_8 hold53 (.A(net379),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\funct3_s2[2] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net370),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_002_),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_004_),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net350),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\data_reg[13] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\funct3_s2[0] ),
    .X(net397));
 sky130_fd_sc_hd__buf_4 hold63 (.A(\data_reg[10] ),
    .X(net392));
 sky130_fd_sc_hd__buf_8 hold65 (.A(net362),
    .X(net399));
 sky130_fd_sc_hd__buf_8 hold68 (.A(\data_reg[29] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net352),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_4 hold72 (.A(net438),
    .X(net401));
 sky130_fd_sc_hd__buf_6 hold8 (.A(net354),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net392),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\data_reg[31] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\data_reg[16] ),
    .X(net418));
 sky130_fd_sc_hd__buf_4 hold9 (.A(net466),
    .X(net338));
 sky130_fd_sc_hd__buf_4 hold94 (.A(\data_reg[17] ),
    .X(net423));
 sky130_fd_sc_hd__buf_8 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_16 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(io_in[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_8 input5 (.A(io_in[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 max_cap107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 max_cap115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 max_cap121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 max_cap127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__buf_2 max_cap151 (.A(net152),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 max_cap172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__buf_2 max_cap177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 max_cap18 (.A(net344),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 max_cap203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 max_cap224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 max_cap27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 max_cap271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_2 max_cap279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_2 max_cap280 (.A(net281),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_2 max_cap285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 max_cap289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__buf_2 max_cap33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 max_cap40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 max_cap47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 max_cap53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 max_cap58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 max_cap68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 max_cap78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 max_cap83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 max_cap99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__conb_1 osiris_i_mem_316 (.LO(net316));
 sky130_fd_sc_hd__conb_1 osiris_i_mem_317 (.LO(net317));
 sky130_fd_sc_hd__conb_1 osiris_i_mem_318 (.LO(net318));
 sky130_fd_sc_hd__conb_1 osiris_i_mem_319 (.LO(net319));
 sky130_fd_sc_hd__conb_1 osiris_i_mem_320 (.LO(net320));
 sky130_fd_sc_hd__conb_1 osiris_i_mem_321 (.LO(net321));
 sky130_fd_sc_hd__conb_1 osiris_i_mem_322 (.LO(net322));
 sky130_fd_sc_hd__buf_12 output6 (.A(net6),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_12 output7 (.A(net7),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_1 wire1 (.A(net9),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 wire10 (.A(\mux_funct3[1] ),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 wire100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__buf_2 wire101 (.A(\core_instr_ID[21] ),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 wire102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__buf_2 wire103 (.A(\core_instr_ID[20] ),
    .X(net103));
 sky130_fd_sc_hd__buf_1 wire104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__buf_4 wire105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 wire106 (.A(net108),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 wire108 (.A(\core_instr_ID[1] ),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 wire109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 wire11 (.A(\mux_funct3[0] ),
    .X(net11));
 sky130_fd_sc_hd__buf_2 wire110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 wire111 (.A(\core_instr_ID[19] ),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 wire112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 wire113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 wire114 (.A(net116),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 wire116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__buf_2 wire117 (.A(\core_instr_ID[18] ),
    .X(net117));
 sky130_fd_sc_hd__buf_4 wire118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 wire119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 wire120 (.A(net122),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 wire122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 wire123 (.A(\core_instr_ID[17] ),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 wire124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 wire125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__buf_2 wire126 (.A(\core_instr_ID[16] ),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 wire128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__buf_2 wire129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 wire130 (.A(\core_instr_ID[15] ),
    .X(net130));
 sky130_fd_sc_hd__buf_2 wire131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 wire132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__buf_2 wire133 (.A(\core_instr_ID[14] ),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 wire134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_2 wire135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 wire136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__buf_2 wire137 (.A(\core_instr_ID[13] ),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_2 wire138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 wire139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 wire140 (.A(net141),
    .X(net140));
 sky130_fd_sc_hd__buf_2 wire141 (.A(\core_instr_ID[12] ),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 wire142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__buf_8 wire143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 wire144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 wire145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_2 wire146 (.A(\core_instr_ID[11] ),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 wire147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__buf_2 wire148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__buf_2 wire149 (.A(\core_instr_ID[10] ),
    .X(net149));
 sky130_fd_sc_hd__buf_2 wire150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_2 wire152 (.A(\core_instr_ID[0] ),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 wire153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 wire154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 wire155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 wire156 (.A(\core_read_data_M[9] ),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 wire157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 wire158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 wire159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 wire160 (.A(\core_read_data_M[8] ),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 wire161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 wire162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 wire163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 wire164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 wire165 (.A(\core_read_data_M[7] ),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 wire166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__buf_2 wire167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 wire168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__buf_2 wire169 (.A(\core_read_data_M[6] ),
    .X(net169));
 sky130_fd_sc_hd__buf_8 wire170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__buf_1 wire171 (.A(net173),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 wire173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 wire174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__buf_2 wire175 (.A(\core_read_data_M[5] ),
    .X(net175));
 sky130_fd_sc_hd__buf_2 wire176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__buf_6 wire178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 wire179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 wire180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__buf_2 wire181 (.A(\core_read_data_M[4] ),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 wire182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__buf_6 wire183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_2 wire184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 wire185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 wire186 (.A(\core_read_data_M[3] ),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_2 wire187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__buf_6 wire188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__buf_6 wire189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 wire190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__buf_8 wire191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 wire192 (.A(\core_read_data_M[31] ),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_2 wire193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__buf_6 wire194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__buf_6 wire195 (.A(net196),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 wire196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_4 wire197 (.A(net198),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 wire198 (.A(\core_read_data_M[30] ),
    .X(net198));
 sky130_fd_sc_hd__buf_6 wire199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_1 wire2 (.A(net8),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 wire200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 wire201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 wire202 (.A(net384),
    .X(net202));
 sky130_fd_sc_hd__buf_6 wire204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__buf_4 wire205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__buf_6 wire206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 wire207 (.A(\core_read_data_M[29] ),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 wire208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__buf_6 wire209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__buf_6 wire210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 wire211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__buf_8 wire212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 wire213 (.A(\core_read_data_M[28] ),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 wire214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_6 wire215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__buf_1 wire216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_4 wire217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_2 wire218 (.A(\core_read_data_M[27] ),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 wire219 (.A(net220),
    .X(net219));
 sky130_fd_sc_hd__buf_6 wire220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_2 wire221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 wire222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 wire223 (.A(\core_read_data_M[26] ),
    .X(net223));
 sky130_fd_sc_hd__buf_6 wire225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__buf_6 wire226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 wire227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 wire228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__buf_8 wire229 (.A(\core_read_data_M[25] ),
    .X(net229));
 sky130_fd_sc_hd__buf_2 wire23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 wire230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__buf_6 wire231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 wire232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_4 wire233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 wire234 (.A(\core_read_data_M[24] ),
    .X(net234));
 sky130_fd_sc_hd__buf_4 wire235 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__buf_6 wire236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__buf_6 wire237 (.A(net238),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 wire238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__buf_4 wire239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__buf_2 wire24 (.A(\core_instr_ID[9] ),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 wire240 (.A(\core_read_data_M[23] ),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 wire241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__buf_6 wire242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 wire243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_2 wire244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__buf_6 wire245 (.A(\core_read_data_M[22] ),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_2 wire246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__buf_6 wire247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 wire248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 wire249 (.A(net250),
    .X(net249));
 sky130_fd_sc_hd__buf_1 wire25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 wire250 (.A(\core_read_data_M[21] ),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 wire251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__buf_6 wire252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 wire253 (.A(net254),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_4 wire254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 wire255 (.A(\core_read_data_M[20] ),
    .X(net255));
 sky130_fd_sc_hd__buf_4 wire256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_2 wire257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 wire258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 wire259 (.A(\core_read_data_M[1] ),
    .X(net259));
 sky130_fd_sc_hd__buf_6 wire26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_6 wire260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__buf_6 wire261 (.A(net262),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 wire262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 wire263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__buf_6 wire264 (.A(\core_read_data_M[19] ),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_2 wire265 (.A(net266),
    .X(net265));
 sky130_fd_sc_hd__buf_6 wire266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_2 wire267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_4 wire268 (.A(net269),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_2 wire269 (.A(\core_read_data_M[18] ),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_2 wire270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_2 wire272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_4 wire273 (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_2 wire274 (.A(\core_read_data_M[17] ),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_2 wire275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_2 wire276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_2 wire277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 wire278 (.A(\core_read_data_M[16] ),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_2 wire28 (.A(\core_instr_ID[8] ),
    .X(net28));
 sky130_fd_sc_hd__buf_6 wire281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_2 wire282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 wire283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_2 wire284 (.A(\core_read_data_M[15] ),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_2 wire286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 wire287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 wire288 (.A(\core_read_data_M[14] ),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_2 wire29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 wire290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_2 wire291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_4 wire292 (.A(\core_read_data_M[13] ),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_2 wire293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_2 wire294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_2 wire295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 wire296 (.A(\core_read_data_M[12] ),
    .X(net296));
 sky130_fd_sc_hd__buf_6 wire297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_2 wire298 (.A(net299),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_2 wire299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__buf_1 wire3 (.A(net10),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_2 wire30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 wire300 (.A(\core_read_data_M[11] ),
    .X(net300));
 sky130_fd_sc_hd__buf_6 wire301 (.A(net302),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_2 wire302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 wire303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_4 wire304 (.A(\core_read_data_M[10] ),
    .X(net304));
 sky130_fd_sc_hd__buf_6 wire305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_2 wire306 (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_2 wire307 (.A(net308),
    .X(net307));
 sky130_fd_sc_hd__buf_2 wire308 (.A(\core_read_data_M[0] ),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_2 wire31 (.A(\core_instr_ID[7] ),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 wire32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__buf_2 wire34 (.A(\core_instr_ID[6] ),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 wire35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 wire36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 wire37 (.A(\core_instr_ID[5] ),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 wire38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_8 wire39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__buf_1 wire4 (.A(net11),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_2 wire41 (.A(\core_instr_ID[4] ),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 wire42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__buf_2 wire43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 wire44 (.A(\core_instr_ID[3] ),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 wire45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_8 wire46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 wire48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 wire49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__buf_2 wire5 (.A(\core_read_data_M[2] ),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_2 wire50 (.A(\core_instr_ID[31] ),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 wire51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 wire52 (.A(net54),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 wire54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 wire55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 wire56 (.A(\core_instr_ID[30] ),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 wire57 (.A(net59),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 wire59 (.A(\core_instr_ID[2] ),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 wire60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 wire61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 wire62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 wire63 (.A(\core_instr_ID[29] ),
    .X(net63));
 sky130_fd_sc_hd__buf_6 wire64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 wire65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__buf_6 wire66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 wire67 (.A(net69),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 wire69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 wire70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 wire71 (.A(\core_instr_ID[28] ),
    .X(net71));
 sky130_fd_sc_hd__buf_4 wire72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__buf_2 wire73 (.A(net74),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 wire74 (.A(\core_instr_ID[27] ),
    .X(net74));
 sky130_fd_sc_hd__buf_4 wire75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 wire76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 wire77 (.A(net79),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 wire79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 wire8 (.A(\mux_funct3[3] ),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 wire80 (.A(\core_instr_ID[26] ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 wire81 (.A(net82),
    .X(net81));
 sky130_fd_sc_hd__buf_8 wire82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 wire84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 wire85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 wire86 (.A(\core_instr_ID[25] ),
    .X(net86));
 sky130_fd_sc_hd__buf_2 wire87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 wire88 (.A(net89),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 wire89 (.A(\core_instr_ID[24] ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 wire9 (.A(\mux_funct3[2] ),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 wire90 (.A(net92),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 wire91 (.A(net92),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 wire92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 wire93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 wire94 (.A(\core_instr_ID[23] ),
    .X(net94));
 sky130_fd_sc_hd__buf_4 wire95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__buf_2 wire96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 wire97 (.A(\core_instr_ID[22] ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 wire98 (.A(net99),
    .X(net98));
 assign io_oeb[0] = net316;
 assign io_oeb[1] = net317;
 assign io_oeb[2] = net318;
 assign io_oeb[3] = net319;
 assign io_oeb[4] = net320;
 assign io_oeb[5] = net321;
 assign io_oeb[6] = net322;
endmodule

