magic
tech sky130A
magscale 1 2
timestamp 1730780735
<< obsli1 >>
rect 2760 2703 97152 97393
<< obsm1 >>
rect 14 2672 98610 97424
<< metal2 >>
rect 3882 99200 3938 100000
rect 9034 99200 9090 100000
rect 14186 99200 14242 100000
rect 19338 99200 19394 100000
rect 24490 99200 24546 100000
rect 29642 99200 29698 100000
rect 34794 99200 34850 100000
rect 40590 99200 40646 100000
rect 45742 99200 45798 100000
rect 50894 99200 50950 100000
rect 56046 99200 56102 100000
rect 61198 99200 61254 100000
rect 66350 99200 66406 100000
rect 71502 99200 71558 100000
rect 76654 99200 76710 100000
rect 81806 99200 81862 100000
rect 86958 99200 87014 100000
rect 92110 99200 92166 100000
rect 97262 99200 97318 100000
rect 18 0 74 800
rect 5170 0 5226 800
rect 10322 0 10378 800
rect 15474 0 15530 800
rect 20626 0 20682 800
rect 25778 0 25834 800
rect 30930 0 30986 800
rect 36082 0 36138 800
rect 41234 0 41290 800
rect 46386 0 46442 800
rect 51538 0 51594 800
rect 56690 0 56746 800
rect 61842 0 61898 800
rect 67638 0 67694 800
rect 72790 0 72846 800
rect 77942 0 77998 800
rect 83094 0 83150 800
rect 88246 0 88302 800
rect 93398 0 93454 800
rect 98550 0 98606 800
<< obsm2 >>
rect 20 99144 3826 99362
rect 3994 99144 8978 99362
rect 9146 99144 14130 99362
rect 14298 99144 19282 99362
rect 19450 99144 24434 99362
rect 24602 99144 29586 99362
rect 29754 99144 34738 99362
rect 34906 99144 40534 99362
rect 40702 99144 45686 99362
rect 45854 99144 50838 99362
rect 51006 99144 55990 99362
rect 56158 99144 61142 99362
rect 61310 99144 66294 99362
rect 66462 99144 71446 99362
rect 71614 99144 76598 99362
rect 76766 99144 81750 99362
rect 81918 99144 86902 99362
rect 87070 99144 92054 99362
rect 92222 99144 97206 99362
rect 97374 99144 98604 99362
rect 20 856 98604 99144
rect 130 800 5114 856
rect 5282 800 10266 856
rect 10434 800 15418 856
rect 15586 800 20570 856
rect 20738 800 25722 856
rect 25890 800 30874 856
rect 31042 800 36026 856
rect 36194 800 41178 856
rect 41346 800 46330 856
rect 46498 800 51482 856
rect 51650 800 56634 856
rect 56802 800 61786 856
rect 61954 800 67582 856
rect 67750 800 72734 856
rect 72902 800 77886 856
rect 78054 800 83038 856
rect 83206 800 88190 856
rect 88358 800 93342 856
rect 93510 800 98494 856
<< metal3 >>
rect 0 98608 800 98728
rect 99200 96568 100000 96688
rect 0 93168 800 93288
rect 99200 91128 100000 91248
rect 0 87728 800 87848
rect 99200 85688 100000 85808
rect 0 82288 800 82408
rect 99200 80248 100000 80368
rect 0 76848 800 76968
rect 99200 74808 100000 74928
rect 0 71408 800 71528
rect 99200 69368 100000 69488
rect 0 65288 800 65408
rect 99200 63928 100000 64048
rect 0 59848 800 59968
rect 99200 58488 100000 58608
rect 0 54408 800 54528
rect 99200 53048 100000 53168
rect 0 48968 800 49088
rect 99200 47608 100000 47728
rect 0 43528 800 43648
rect 99200 42168 100000 42288
rect 0 38088 800 38208
rect 99200 36728 100000 36848
rect 0 32648 800 32768
rect 99200 31288 100000 31408
rect 0 27208 800 27328
rect 99200 25168 100000 25288
rect 0 21768 800 21888
rect 99200 19728 100000 19848
rect 0 16328 800 16448
rect 99200 14288 100000 14408
rect 0 10888 800 11008
rect 99200 8848 100000 8968
rect 0 5448 800 5568
rect 99200 3408 100000 3528
<< obsm3 >>
rect 880 98528 99200 98701
rect 800 96768 99200 98528
rect 800 96488 99120 96768
rect 800 93368 99200 96488
rect 880 93088 99200 93368
rect 800 91328 99200 93088
rect 800 91048 99120 91328
rect 800 87928 99200 91048
rect 880 87648 99200 87928
rect 800 85888 99200 87648
rect 800 85608 99120 85888
rect 800 82488 99200 85608
rect 880 82208 99200 82488
rect 800 80448 99200 82208
rect 800 80168 99120 80448
rect 800 77048 99200 80168
rect 880 76768 99200 77048
rect 800 75008 99200 76768
rect 800 74728 99120 75008
rect 800 71608 99200 74728
rect 880 71328 99200 71608
rect 800 69568 99200 71328
rect 800 69288 99120 69568
rect 800 65488 99200 69288
rect 880 65208 99200 65488
rect 800 64128 99200 65208
rect 800 63848 99120 64128
rect 800 60048 99200 63848
rect 880 59768 99200 60048
rect 800 58688 99200 59768
rect 800 58408 99120 58688
rect 800 54608 99200 58408
rect 880 54328 99200 54608
rect 800 53248 99200 54328
rect 800 52968 99120 53248
rect 800 49168 99200 52968
rect 880 48888 99200 49168
rect 800 47808 99200 48888
rect 800 47528 99120 47808
rect 800 43728 99200 47528
rect 880 43448 99200 43728
rect 800 42368 99200 43448
rect 800 42088 99120 42368
rect 800 38288 99200 42088
rect 880 38008 99200 38288
rect 800 36928 99200 38008
rect 800 36648 99120 36928
rect 800 32848 99200 36648
rect 880 32568 99200 32848
rect 800 31488 99200 32568
rect 800 31208 99120 31488
rect 800 27408 99200 31208
rect 880 27128 99200 27408
rect 800 25368 99200 27128
rect 800 25088 99120 25368
rect 800 21968 99200 25088
rect 880 21688 99200 21968
rect 800 19928 99200 21688
rect 800 19648 99120 19928
rect 800 16528 99200 19648
rect 880 16248 99200 16528
rect 800 14488 99200 16248
rect 800 14208 99120 14488
rect 800 11088 99200 14208
rect 880 10808 99200 11088
rect 800 9048 99200 10808
rect 800 8768 99120 9048
rect 800 5648 99200 8768
rect 880 5368 99200 5648
rect 800 3608 99200 5368
rect 800 3328 99120 3608
rect 800 2687 99200 3328
<< metal4 >>
rect 5864 2672 6184 97424
rect 6524 2672 6844 97424
rect 41864 2672 42184 97424
rect 42524 2672 42844 97424
rect 77864 2672 78184 97424
rect 78524 2672 78844 97424
<< obsm4 >>
rect 25819 3027 41784 96933
rect 42264 3027 42444 96933
rect 42924 3027 77784 96933
rect 78264 3027 78444 96933
rect 78924 3027 95621 96933
<< labels >>
rlabel metal3 s 0 10888 800 11008 6 clk
port 1 nsew signal input
rlabel metal3 s 99200 36728 100000 36848 6 rst
port 2 nsew signal input
rlabel metal4 s 5864 2672 6184 97424 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 41864 2672 42184 97424 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 77864 2672 78184 97424 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 6524 2672 6844 97424 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 42524 2672 42844 97424 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 78524 2672 78844 97424 6 vssd1
port 4 nsew ground bidirectional
rlabel metal2 s 77942 0 77998 800 6 wb_ack_o
port 5 nsew signal output
rlabel metal3 s 99200 63928 100000 64048 6 wb_adr_i[0]
port 6 nsew signal input
rlabel metal3 s 99200 14288 100000 14408 6 wb_adr_i[1]
port 7 nsew signal input
rlabel metal2 s 19338 99200 19394 100000 6 wb_adr_i[2]
port 8 nsew signal input
rlabel metal2 s 71502 99200 71558 100000 6 wb_adr_i[3]
port 9 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wb_adr_i[4]
port 10 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 wb_cyc_i
port 11 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 wb_dat_i[0]
port 12 nsew signal input
rlabel metal2 s 97262 99200 97318 100000 6 wb_dat_i[10]
port 13 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wb_dat_i[11]
port 14 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 wb_dat_i[12]
port 15 nsew signal input
rlabel metal3 s 99200 19728 100000 19848 6 wb_dat_i[13]
port 16 nsew signal input
rlabel metal3 s 99200 58488 100000 58608 6 wb_dat_i[14]
port 17 nsew signal input
rlabel metal3 s 99200 74808 100000 74928 6 wb_dat_i[15]
port 18 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 wb_dat_i[16]
port 19 nsew signal input
rlabel metal3 s 99200 80248 100000 80368 6 wb_dat_i[17]
port 20 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 wb_dat_i[18]
port 21 nsew signal input
rlabel metal3 s 99200 25168 100000 25288 6 wb_dat_i[19]
port 22 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 wb_dat_i[1]
port 23 nsew signal input
rlabel metal2 s 66350 99200 66406 100000 6 wb_dat_i[20]
port 24 nsew signal input
rlabel metal3 s 99200 69368 100000 69488 6 wb_dat_i[21]
port 25 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 wb_dat_i[22]
port 26 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 wb_dat_i[23]
port 27 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wb_dat_i[24]
port 28 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wb_dat_i[25]
port 29 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 wb_dat_i[26]
port 30 nsew signal input
rlabel metal2 s 9034 99200 9090 100000 6 wb_dat_i[27]
port 31 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 wb_dat_i[28]
port 32 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 wb_dat_i[29]
port 33 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 wb_dat_i[2]
port 34 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wb_dat_i[30]
port 35 nsew signal input
rlabel metal2 s 34794 99200 34850 100000 6 wb_dat_i[31]
port 36 nsew signal input
rlabel metal2 s 3882 99200 3938 100000 6 wb_dat_i[3]
port 37 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 wb_dat_i[4]
port 38 nsew signal input
rlabel metal2 s 45742 99200 45798 100000 6 wb_dat_i[5]
port 39 nsew signal input
rlabel metal2 s 92110 99200 92166 100000 6 wb_dat_i[6]
port 40 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 wb_dat_i[7]
port 41 nsew signal input
rlabel metal2 s 50894 99200 50950 100000 6 wb_dat_i[8]
port 42 nsew signal input
rlabel metal3 s 99200 8848 100000 8968 6 wb_dat_i[9]
port 43 nsew signal input
rlabel metal3 s 99200 31288 100000 31408 6 wb_dat_o[0]
port 44 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 wb_dat_o[10]
port 45 nsew signal output
rlabel metal3 s 99200 42168 100000 42288 6 wb_dat_o[11]
port 46 nsew signal output
rlabel metal2 s 40590 99200 40646 100000 6 wb_dat_o[12]
port 47 nsew signal output
rlabel metal2 s 61198 99200 61254 100000 6 wb_dat_o[13]
port 48 nsew signal output
rlabel metal3 s 0 98608 800 98728 6 wb_dat_o[14]
port 49 nsew signal output
rlabel metal2 s 18 0 74 800 6 wb_dat_o[15]
port 50 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 wb_dat_o[16]
port 51 nsew signal output
rlabel metal2 s 56046 99200 56102 100000 6 wb_dat_o[17]
port 52 nsew signal output
rlabel metal2 s 76654 99200 76710 100000 6 wb_dat_o[18]
port 53 nsew signal output
rlabel metal3 s 99200 96568 100000 96688 6 wb_dat_o[19]
port 54 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 wb_dat_o[1]
port 55 nsew signal output
rlabel metal3 s 0 71408 800 71528 6 wb_dat_o[20]
port 56 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 wb_dat_o[21]
port 57 nsew signal output
rlabel metal3 s 99200 91128 100000 91248 6 wb_dat_o[22]
port 58 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 wb_dat_o[23]
port 59 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 wb_dat_o[24]
port 60 nsew signal output
rlabel metal3 s 99200 85688 100000 85808 6 wb_dat_o[25]
port 61 nsew signal output
rlabel metal3 s 99200 3408 100000 3528 6 wb_dat_o[26]
port 62 nsew signal output
rlabel metal2 s 24490 99200 24546 100000 6 wb_dat_o[27]
port 63 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 wb_dat_o[28]
port 64 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wb_dat_o[29]
port 65 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 wb_dat_o[2]
port 66 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 wb_dat_o[30]
port 67 nsew signal output
rlabel metal3 s 99200 53048 100000 53168 6 wb_dat_o[31]
port 68 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 wb_dat_o[3]
port 69 nsew signal output
rlabel metal2 s 86958 99200 87014 100000 6 wb_dat_o[4]
port 70 nsew signal output
rlabel metal2 s 81806 99200 81862 100000 6 wb_dat_o[5]
port 71 nsew signal output
rlabel metal2 s 14186 99200 14242 100000 6 wb_dat_o[6]
port 72 nsew signal output
rlabel metal2 s 29642 99200 29698 100000 6 wb_dat_o[7]
port 73 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 wb_dat_o[8]
port 74 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 wb_dat_o[9]
port 75 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 wb_stb_i
port 76 nsew signal input
rlabel metal3 s 99200 47608 100000 47728 6 wb_we_i
port 77 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17884574
string GDS_FILE /home/roliveira/Desktop/osiris_i/openlane/mem/runs/metal/results/signoff/mem.magic.gds
string GDS_START 390084
<< end >>

