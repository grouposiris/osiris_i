VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.210 BY 397.090 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END clk
  PIN i_instr_ID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 393.090 196.790 397.090 ;
    END
  END i_instr_ID[0]
  PIN i_instr_ID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 380.840 400.210 381.440 ;
    END
  END i_instr_ID[10]
  PIN i_instr_ID[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 319.640 400.210 320.240 ;
    END
  END i_instr_ID[11]
  PIN i_instr_ID[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 235.150 393.090 235.430 397.090 ;
    END
  END i_instr_ID[12]
  PIN i_instr_ID[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END i_instr_ID[13]
  PIN i_instr_ID[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 357.510 393.090 357.790 397.090 ;
    END
  END i_instr_ID[14]
  PIN i_instr_ID[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END i_instr_ID[15]
  PIN i_instr_ID[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 6.840 400.210 7.440 ;
    END
  END i_instr_ID[16]
  PIN i_instr_ID[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 244.810 393.090 245.090 397.090 ;
    END
  END i_instr_ID[17]
  PIN i_instr_ID[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 108.840 400.210 109.440 ;
    END
  END i_instr_ID[18]
  PIN i_instr_ID[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 221.040 400.210 221.640 ;
    END
  END i_instr_ID[19]
  PIN i_instr_ID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 393.090 138.830 397.090 ;
    END
  END i_instr_ID[1]
  PIN i_instr_ID[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END i_instr_ID[20]
  PIN i_instr_ID[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 393.090 177.470 397.090 ;
    END
  END i_instr_ID[21]
  PIN i_instr_ID[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END i_instr_ID[22]
  PIN i_instr_ID[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END i_instr_ID[23]
  PIN i_instr_ID[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END i_instr_ID[24]
  PIN i_instr_ID[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 180.240 400.210 180.840 ;
    END
  END i_instr_ID[25]
  PIN i_instr_ID[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 393.090 42.230 397.090 ;
    END
  END i_instr_ID[26]
  PIN i_instr_ID[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 270.570 393.090 270.850 397.090 ;
    END
  END i_instr_ID[27]
  PIN i_instr_ID[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END i_instr_ID[28]
  PIN i_instr_ID[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END i_instr_ID[29]
  PIN i_instr_ID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 396.150 393.090 396.430 397.090 ;
    END
  END i_instr_ID[2]
  PIN i_instr_ID[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END i_instr_ID[30]
  PIN i_instr_ID[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END i_instr_ID[31]
  PIN i_instr_ID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 37.440 400.210 38.040 ;
    END
  END i_instr_ID[3]
  PIN i_instr_ID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END i_instr_ID[4]
  PIN i_instr_ID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END i_instr_ID[5]
  PIN i_instr_ID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END i_instr_ID[6]
  PIN i_instr_ID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END i_instr_ID[7]
  PIN i_instr_ID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 393.090 109.850 397.090 ;
    END
  END i_instr_ID[8]
  PIN i_instr_ID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 225.490 393.090 225.770 397.090 ;
    END
  END i_instr_ID[9]
  PIN i_read_data_M[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 367.170 393.090 367.450 397.090 ;
    END
  END i_read_data_M[0]
  PIN i_read_data_M[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END i_read_data_M[10]
  PIN i_read_data_M[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 393.090 51.890 397.090 ;
    END
  END i_read_data_M[11]
  PIN i_read_data_M[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 309.440 400.210 310.040 ;
    END
  END i_read_data_M[12]
  PIN i_read_data_M[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 386.490 393.090 386.770 397.090 ;
    END
  END i_read_data_M[13]
  PIN i_read_data_M[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 289.040 400.210 289.640 ;
    END
  END i_read_data_M[14]
  PIN i_read_data_M[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END i_read_data_M[15]
  PIN i_read_data_M[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END i_read_data_M[16]
  PIN i_read_data_M[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END i_read_data_M[17]
  PIN i_read_data_M[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 159.840 400.210 160.440 ;
    END
  END i_read_data_M[18]
  PIN i_read_data_M[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END i_read_data_M[19]
  PIN i_read_data_M[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END i_read_data_M[1]
  PIN i_read_data_M[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 17.040 400.210 17.640 ;
    END
  END i_read_data_M[20]
  PIN i_read_data_M[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 157.870 393.090 158.150 397.090 ;
    END
  END i_read_data_M[21]
  PIN i_read_data_M[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END i_read_data_M[22]
  PIN i_read_data_M[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END i_read_data_M[23]
  PIN i_read_data_M[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END i_read_data_M[24]
  PIN i_read_data_M[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 186.850 393.090 187.130 397.090 ;
    END
  END i_read_data_M[25]
  PIN i_read_data_M[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 393.090 32.570 397.090 ;
    END
  END i_read_data_M[26]
  PIN i_read_data_M[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 299.240 400.210 299.840 ;
    END
  END i_read_data_M[27]
  PIN i_read_data_M[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END i_read_data_M[28]
  PIN i_read_data_M[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END i_read_data_M[29]
  PIN i_read_data_M[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 148.210 393.090 148.490 397.090 ;
    END
  END i_read_data_M[2]
  PIN i_read_data_M[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 88.440 400.210 89.040 ;
    END
  END i_read_data_M[30]
  PIN i_read_data_M[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 340.040 400.210 340.640 ;
    END
  END i_read_data_M[31]
  PIN i_read_data_M[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 129.240 400.210 129.840 ;
    END
  END i_read_data_M[3]
  PIN i_read_data_M[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END i_read_data_M[4]
  PIN i_read_data_M[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 47.640 400.210 48.240 ;
    END
  END i_read_data_M[5]
  PIN i_read_data_M[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END i_read_data_M[6]
  PIN i_read_data_M[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END i_read_data_M[7]
  PIN i_read_data_M[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.210 360.440 400.210 361.040 ;
    END
  END i_read_data_M[8]
  PIN i_read_data_M[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END i_read_data_M[9]
  PIN o_data_addr_M[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 376.830 393.090 377.110 397.090 ;
    END
  END o_data_addr_M[0]
  PIN o_data_addr_M[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END o_data_addr_M[10]
  PIN o_data_addr_M[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END o_data_addr_M[11]
  PIN o_data_addr_M[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 280.230 393.090 280.510 397.090 ;
    END
  END o_data_addr_M[12]
  PIN o_data_addr_M[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 260.910 393.090 261.190 397.090 ;
    END
  END o_data_addr_M[13]
  PIN o_data_addr_M[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 393.090 129.170 397.090 ;
    END
  END o_data_addr_M[14]
  PIN o_data_addr_M[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END o_data_addr_M[15]
  PIN o_data_addr_M[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 22.630 393.090 22.910 397.090 ;
    END
  END o_data_addr_M[16]
  PIN o_data_addr_M[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 350.240 400.210 350.840 ;
    END
  END o_data_addr_M[17]
  PIN o_data_addr_M[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END o_data_addr_M[18]
  PIN o_data_addr_M[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END o_data_addr_M[19]
  PIN o_data_addr_M[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 278.840 400.210 279.440 ;
    END
  END o_data_addr_M[1]
  PIN o_data_addr_M[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END o_data_addr_M[20]
  PIN o_data_addr_M[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END o_data_addr_M[21]
  PIN o_data_addr_M[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 238.040 400.210 238.640 ;
    END
  END o_data_addr_M[22]
  PIN o_data_addr_M[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END o_data_addr_M[23]
  PIN o_data_addr_M[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 78.240 400.210 78.840 ;
    END
  END o_data_addr_M[24]
  PIN o_data_addr_M[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 393.090 100.190 397.090 ;
    END
  END o_data_addr_M[25]
  PIN o_data_addr_M[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 149.640 400.210 150.240 ;
    END
  END o_data_addr_M[26]
  PIN o_data_addr_M[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END o_data_addr_M[27]
  PIN o_data_addr_M[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 347.850 393.090 348.130 397.090 ;
    END
  END o_data_addr_M[28]
  PIN o_data_addr_M[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 170.040 400.210 170.640 ;
    END
  END o_data_addr_M[29]
  PIN o_data_addr_M[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END o_data_addr_M[2]
  PIN o_data_addr_M[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END o_data_addr_M[30]
  PIN o_data_addr_M[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 251.250 393.090 251.530 397.090 ;
    END
  END o_data_addr_M[31]
  PIN o_data_addr_M[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END o_data_addr_M[3]
  PIN o_data_addr_M[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END o_data_addr_M[4]
  PIN o_data_addr_M[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 12.970 393.090 13.250 397.090 ;
    END
  END o_data_addr_M[5]
  PIN o_data_addr_M[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 61.270 393.090 61.550 397.090 ;
    END
  END o_data_addr_M[6]
  PIN o_data_addr_M[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 309.210 393.090 309.490 397.090 ;
    END
  END o_data_addr_M[7]
  PIN o_data_addr_M[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 318.870 393.090 319.150 397.090 ;
    END
  END o_data_addr_M[8]
  PIN o_data_addr_M[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 299.550 393.090 299.830 397.090 ;
    END
  END o_data_addr_M[9]
  PIN o_mem_write_M
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END o_mem_write_M
  PIN o_pc_IF[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END o_pc_IF[0]
  PIN o_pc_IF[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 27.240 400.210 27.840 ;
    END
  END o_pc_IF[10]
  PIN o_pc_IF[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END o_pc_IF[11]
  PIN o_pc_IF[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 119.230 393.090 119.510 397.090 ;
    END
  END o_pc_IF[12]
  PIN o_pc_IF[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 200.640 400.210 201.240 ;
    END
  END o_pc_IF[13]
  PIN o_pc_IF[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 328.530 393.090 328.810 397.090 ;
    END
  END o_pc_IF[14]
  PIN o_pc_IF[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END o_pc_IF[15]
  PIN o_pc_IF[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END o_pc_IF[16]
  PIN o_pc_IF[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 210.840 400.210 211.440 ;
    END
  END o_pc_IF[17]
  PIN o_pc_IF[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 167.530 393.090 167.810 397.090 ;
    END
  END o_pc_IF[18]
  PIN o_pc_IF[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 139.440 400.210 140.040 ;
    END
  END o_pc_IF[19]
  PIN o_pc_IF[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END o_pc_IF[1]
  PIN o_pc_IF[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END o_pc_IF[20]
  PIN o_pc_IF[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 268.640 400.210 269.240 ;
    END
  END o_pc_IF[21]
  PIN o_pc_IF[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END o_pc_IF[22]
  PIN o_pc_IF[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END o_pc_IF[23]
  PIN o_pc_IF[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 98.640 400.210 99.240 ;
    END
  END o_pc_IF[24]
  PIN o_pc_IF[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END o_pc_IF[25]
  PIN o_pc_IF[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END o_pc_IF[26]
  PIN o_pc_IF[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 393.090 90.530 397.090 ;
    END
  END o_pc_IF[27]
  PIN o_pc_IF[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END o_pc_IF[28]
  PIN o_pc_IF[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END o_pc_IF[29]
  PIN o_pc_IF[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END o_pc_IF[2]
  PIN o_pc_IF[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 57.840 400.210 58.440 ;
    END
  END o_pc_IF[30]
  PIN o_pc_IF[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 329.840 400.210 330.440 ;
    END
  END o_pc_IF[31]
  PIN o_pc_IF[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 231.240 400.210 231.840 ;
    END
  END o_pc_IF[3]
  PIN o_pc_IF[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END o_pc_IF[4]
  PIN o_pc_IF[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END o_pc_IF[5]
  PIN o_pc_IF[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 119.040 400.210 119.640 ;
    END
  END o_pc_IF[6]
  PIN o_pc_IF[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END o_pc_IF[7]
  PIN o_pc_IF[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 248.240 400.210 248.840 ;
    END
  END o_pc_IF[8]
  PIN o_pc_IF[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 370.640 400.210 371.240 ;
    END
  END o_pc_IF[9]
  PIN o_write_data_M[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END o_write_data_M[0]
  PIN o_write_data_M[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 391.040 400.210 391.640 ;
    END
  END o_write_data_M[10]
  PIN o_write_data_M[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END o_write_data_M[11]
  PIN o_write_data_M[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END o_write_data_M[12]
  PIN o_write_data_M[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END o_write_data_M[13]
  PIN o_write_data_M[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END o_write_data_M[14]
  PIN o_write_data_M[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END o_write_data_M[15]
  PIN o_write_data_M[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END o_write_data_M[16]
  PIN o_write_data_M[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 393.090 80.870 397.090 ;
    END
  END o_write_data_M[17]
  PIN o_write_data_M[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 215.830 393.090 216.110 397.090 ;
    END
  END o_write_data_M[18]
  PIN o_write_data_M[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END o_write_data_M[19]
  PIN o_write_data_M[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END o_write_data_M[1]
  PIN o_write_data_M[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END o_write_data_M[20]
  PIN o_write_data_M[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END o_write_data_M[21]
  PIN o_write_data_M[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 206.170 393.090 206.450 397.090 ;
    END
  END o_write_data_M[22]
  PIN o_write_data_M[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END o_write_data_M[23]
  PIN o_write_data_M[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 338.190 393.090 338.470 397.090 ;
    END
  END o_write_data_M[24]
  PIN o_write_data_M[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 68.040 400.210 68.640 ;
    END
  END o_write_data_M[25]
  PIN o_write_data_M[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END o_write_data_M[26]
  PIN o_write_data_M[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END o_write_data_M[27]
  PIN o_write_data_M[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END o_write_data_M[28]
  PIN o_write_data_M[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END o_write_data_M[29]
  PIN o_write_data_M[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END o_write_data_M[2]
  PIN o_write_data_M[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 258.440 400.210 259.040 ;
    END
  END o_write_data_M[30]
  PIN o_write_data_M[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END o_write_data_M[31]
  PIN o_write_data_M[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END o_write_data_M[3]
  PIN o_write_data_M[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 289.890 393.090 290.170 397.090 ;
    END
  END o_write_data_M[4]
  PIN o_write_data_M[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 3.310 393.090 3.590 397.090 ;
    END
  END o_write_data_M[5]
  PIN o_write_data_M[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 393.090 71.210 397.090 ;
    END
  END o_write_data_M[6]
  PIN o_write_data_M[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END o_write_data_M[7]
  PIN o_write_data_M[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END o_write_data_M[8]
  PIN o_write_data_M[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END o_write_data_M[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 396.210 190.440 400.210 191.040 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.320 13.360 30.920 383.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 182.920 13.360 184.520 383.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 336.520 13.360 338.120 383.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 32.620 13.360 34.220 383.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 186.220 13.360 187.820 383.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 339.820 13.360 341.420 383.760 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 13.800 13.515 386.400 383.605 ;
      LAYER met1 ;
        RECT 0.070 11.940 399.670 384.840 ;
      LAYER met2 ;
        RECT 0.100 392.810 3.030 393.450 ;
        RECT 3.870 392.810 12.690 393.450 ;
        RECT 13.530 392.810 22.350 393.450 ;
        RECT 23.190 392.810 32.010 393.450 ;
        RECT 32.850 392.810 41.670 393.450 ;
        RECT 42.510 392.810 51.330 393.450 ;
        RECT 52.170 392.810 60.990 393.450 ;
        RECT 61.830 392.810 70.650 393.450 ;
        RECT 71.490 392.810 80.310 393.450 ;
        RECT 81.150 392.810 89.970 393.450 ;
        RECT 90.810 392.810 99.630 393.450 ;
        RECT 100.470 392.810 109.290 393.450 ;
        RECT 110.130 392.810 118.950 393.450 ;
        RECT 119.790 392.810 128.610 393.450 ;
        RECT 129.450 392.810 138.270 393.450 ;
        RECT 139.110 392.810 147.930 393.450 ;
        RECT 148.770 392.810 157.590 393.450 ;
        RECT 158.430 392.810 167.250 393.450 ;
        RECT 168.090 392.810 176.910 393.450 ;
        RECT 177.750 392.810 186.570 393.450 ;
        RECT 187.410 392.810 196.230 393.450 ;
        RECT 197.070 392.810 205.890 393.450 ;
        RECT 206.730 392.810 215.550 393.450 ;
        RECT 216.390 392.810 225.210 393.450 ;
        RECT 226.050 392.810 234.870 393.450 ;
        RECT 235.710 392.810 244.530 393.450 ;
        RECT 245.370 392.810 250.970 393.450 ;
        RECT 251.810 392.810 260.630 393.450 ;
        RECT 261.470 392.810 270.290 393.450 ;
        RECT 271.130 392.810 279.950 393.450 ;
        RECT 280.790 392.810 289.610 393.450 ;
        RECT 290.450 392.810 299.270 393.450 ;
        RECT 300.110 392.810 308.930 393.450 ;
        RECT 309.770 392.810 318.590 393.450 ;
        RECT 319.430 392.810 328.250 393.450 ;
        RECT 329.090 392.810 337.910 393.450 ;
        RECT 338.750 392.810 347.570 393.450 ;
        RECT 348.410 392.810 357.230 393.450 ;
        RECT 358.070 392.810 366.890 393.450 ;
        RECT 367.730 392.810 376.550 393.450 ;
        RECT 377.390 392.810 386.210 393.450 ;
        RECT 387.050 392.810 395.870 393.450 ;
        RECT 396.710 392.810 399.640 393.450 ;
        RECT 0.100 4.280 399.640 392.810 ;
        RECT 0.650 4.000 6.250 4.280 ;
        RECT 7.090 4.000 15.910 4.280 ;
        RECT 16.750 4.000 25.570 4.280 ;
        RECT 26.410 4.000 35.230 4.280 ;
        RECT 36.070 4.000 44.890 4.280 ;
        RECT 45.730 4.000 54.550 4.280 ;
        RECT 55.390 4.000 64.210 4.280 ;
        RECT 65.050 4.000 73.870 4.280 ;
        RECT 74.710 4.000 83.530 4.280 ;
        RECT 84.370 4.000 93.190 4.280 ;
        RECT 94.030 4.000 102.850 4.280 ;
        RECT 103.690 4.000 112.510 4.280 ;
        RECT 113.350 4.000 122.170 4.280 ;
        RECT 123.010 4.000 131.830 4.280 ;
        RECT 132.670 4.000 141.490 4.280 ;
        RECT 142.330 4.000 151.150 4.280 ;
        RECT 151.990 4.000 160.810 4.280 ;
        RECT 161.650 4.000 170.470 4.280 ;
        RECT 171.310 4.000 180.130 4.280 ;
        RECT 180.970 4.000 189.790 4.280 ;
        RECT 190.630 4.000 199.450 4.280 ;
        RECT 200.290 4.000 209.110 4.280 ;
        RECT 209.950 4.000 218.770 4.280 ;
        RECT 219.610 4.000 228.430 4.280 ;
        RECT 229.270 4.000 238.090 4.280 ;
        RECT 238.930 4.000 247.750 4.280 ;
        RECT 248.590 4.000 257.410 4.280 ;
        RECT 258.250 4.000 267.070 4.280 ;
        RECT 267.910 4.000 276.730 4.280 ;
        RECT 277.570 4.000 286.390 4.280 ;
        RECT 287.230 4.000 296.050 4.280 ;
        RECT 296.890 4.000 305.710 4.280 ;
        RECT 306.550 4.000 312.150 4.280 ;
        RECT 312.990 4.000 321.810 4.280 ;
        RECT 322.650 4.000 331.470 4.280 ;
        RECT 332.310 4.000 341.130 4.280 ;
        RECT 341.970 4.000 350.790 4.280 ;
        RECT 351.630 4.000 360.450 4.280 ;
        RECT 361.290 4.000 370.110 4.280 ;
        RECT 370.950 4.000 379.770 4.280 ;
        RECT 380.610 4.000 389.430 4.280 ;
        RECT 390.270 4.000 399.090 4.280 ;
      LAYER met3 ;
        RECT 4.400 390.640 395.810 391.505 ;
        RECT 4.000 381.840 396.210 390.640 ;
        RECT 4.400 380.440 395.810 381.840 ;
        RECT 4.000 371.640 396.210 380.440 ;
        RECT 4.400 370.240 395.810 371.640 ;
        RECT 4.000 361.440 396.210 370.240 ;
        RECT 4.400 360.040 395.810 361.440 ;
        RECT 4.000 351.240 396.210 360.040 ;
        RECT 4.400 349.840 395.810 351.240 ;
        RECT 4.000 341.040 396.210 349.840 ;
        RECT 4.400 339.640 395.810 341.040 ;
        RECT 4.000 330.840 396.210 339.640 ;
        RECT 4.400 329.440 395.810 330.840 ;
        RECT 4.000 324.040 396.210 329.440 ;
        RECT 4.400 322.640 396.210 324.040 ;
        RECT 4.000 320.640 396.210 322.640 ;
        RECT 4.000 319.240 395.810 320.640 ;
        RECT 4.000 313.840 396.210 319.240 ;
        RECT 4.400 312.440 396.210 313.840 ;
        RECT 4.000 310.440 396.210 312.440 ;
        RECT 4.000 309.040 395.810 310.440 ;
        RECT 4.000 303.640 396.210 309.040 ;
        RECT 4.400 302.240 396.210 303.640 ;
        RECT 4.000 300.240 396.210 302.240 ;
        RECT 4.000 298.840 395.810 300.240 ;
        RECT 4.000 293.440 396.210 298.840 ;
        RECT 4.400 292.040 396.210 293.440 ;
        RECT 4.000 290.040 396.210 292.040 ;
        RECT 4.000 288.640 395.810 290.040 ;
        RECT 4.000 283.240 396.210 288.640 ;
        RECT 4.400 281.840 396.210 283.240 ;
        RECT 4.000 279.840 396.210 281.840 ;
        RECT 4.000 278.440 395.810 279.840 ;
        RECT 4.000 273.040 396.210 278.440 ;
        RECT 4.400 271.640 396.210 273.040 ;
        RECT 4.000 269.640 396.210 271.640 ;
        RECT 4.000 268.240 395.810 269.640 ;
        RECT 4.000 262.840 396.210 268.240 ;
        RECT 4.400 261.440 396.210 262.840 ;
        RECT 4.000 259.440 396.210 261.440 ;
        RECT 4.000 258.040 395.810 259.440 ;
        RECT 4.000 252.640 396.210 258.040 ;
        RECT 4.400 251.240 396.210 252.640 ;
        RECT 4.000 249.240 396.210 251.240 ;
        RECT 4.000 247.840 395.810 249.240 ;
        RECT 4.000 242.440 396.210 247.840 ;
        RECT 4.400 241.040 396.210 242.440 ;
        RECT 4.000 239.040 396.210 241.040 ;
        RECT 4.000 237.640 395.810 239.040 ;
        RECT 4.000 232.240 396.210 237.640 ;
        RECT 4.400 230.840 395.810 232.240 ;
        RECT 4.000 222.040 396.210 230.840 ;
        RECT 4.400 220.640 395.810 222.040 ;
        RECT 4.000 211.840 396.210 220.640 ;
        RECT 4.400 210.440 395.810 211.840 ;
        RECT 4.000 201.640 396.210 210.440 ;
        RECT 4.400 200.240 395.810 201.640 ;
        RECT 4.000 191.440 396.210 200.240 ;
        RECT 4.400 190.040 395.810 191.440 ;
        RECT 4.000 181.240 396.210 190.040 ;
        RECT 4.400 179.840 395.810 181.240 ;
        RECT 4.000 171.040 396.210 179.840 ;
        RECT 4.400 169.640 395.810 171.040 ;
        RECT 4.000 160.840 396.210 169.640 ;
        RECT 4.400 159.440 395.810 160.840 ;
        RECT 4.000 150.640 396.210 159.440 ;
        RECT 4.400 149.240 395.810 150.640 ;
        RECT 4.000 140.440 396.210 149.240 ;
        RECT 4.400 139.040 395.810 140.440 ;
        RECT 4.000 130.240 396.210 139.040 ;
        RECT 4.400 128.840 395.810 130.240 ;
        RECT 4.000 120.040 396.210 128.840 ;
        RECT 4.400 118.640 395.810 120.040 ;
        RECT 4.000 109.840 396.210 118.640 ;
        RECT 4.400 108.440 395.810 109.840 ;
        RECT 4.000 99.640 396.210 108.440 ;
        RECT 4.400 98.240 395.810 99.640 ;
        RECT 4.000 89.440 396.210 98.240 ;
        RECT 4.400 88.040 395.810 89.440 ;
        RECT 4.000 79.240 396.210 88.040 ;
        RECT 4.400 77.840 395.810 79.240 ;
        RECT 4.000 69.040 396.210 77.840 ;
        RECT 4.400 67.640 395.810 69.040 ;
        RECT 4.000 58.840 396.210 67.640 ;
        RECT 4.400 57.440 395.810 58.840 ;
        RECT 4.000 48.640 396.210 57.440 ;
        RECT 4.400 47.240 395.810 48.640 ;
        RECT 4.000 38.440 396.210 47.240 ;
        RECT 4.400 37.040 395.810 38.440 ;
        RECT 4.000 28.240 396.210 37.040 ;
        RECT 4.400 26.840 395.810 28.240 ;
        RECT 4.000 18.040 396.210 26.840 ;
        RECT 4.400 16.640 395.810 18.040 ;
        RECT 4.000 7.840 396.210 16.640 ;
        RECT 4.400 6.975 395.810 7.840 ;
      LAYER met4 ;
        RECT 15.935 15.135 28.920 382.665 ;
        RECT 31.320 15.135 32.220 382.665 ;
        RECT 34.620 15.135 182.520 382.665 ;
        RECT 184.920 15.135 185.820 382.665 ;
        RECT 188.220 15.135 336.120 382.665 ;
        RECT 338.520 15.135 339.420 382.665 ;
        RECT 341.820 15.135 377.825 382.665 ;
  END
END core
END LIBRARY

