VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mem
  CLASS BLOCK ;
  FOREIGN mem ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 183.640 500.000 184.240 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.320 13.360 30.920 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 209.320 13.360 210.920 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 389.320 13.360 390.920 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 32.620 13.360 34.220 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 212.620 13.360 214.220 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 392.620 13.360 394.220 487.120 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 319.640 500.000 320.240 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 71.440 500.000 72.040 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 496.000 96.970 500.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 357.510 496.000 357.790 500.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wb_adr_i[4]
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 486.310 496.000 486.590 500.000 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 98.640 500.000 99.240 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 292.440 500.000 293.040 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 374.040 500.000 374.640 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 401.240 500.000 401.840 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 125.840 500.000 126.440 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 331.750 496.000 332.030 500.000 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 346.840 500.000 347.440 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 496.000 45.450 500.000 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 496.000 174.250 500.000 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 496.000 19.690 500.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 228.710 496.000 228.990 500.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 460.550 496.000 460.830 500.000 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 254.470 496.000 254.750 500.000 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 44.240 500.000 44.840 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 156.440 500.000 157.040 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 210.840 500.000 211.440 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 202.950 496.000 203.230 500.000 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 305.990 496.000 306.270 500.000 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 280.230 496.000 280.510 500.000 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 383.270 496.000 383.550 500.000 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 482.840 500.000 483.440 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 455.640 500.000 456.240 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 428.440 500.000 429.040 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 17.040 500.000 17.640 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 496.000 122.730 500.000 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 265.240 500.000 265.840 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 434.790 496.000 435.070 500.000 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 409.030 496.000 409.310 500.000 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 496.000 71.210 500.000 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 496.000 148.490 500.000 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END wb_dat_o[9]
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 238.040 500.000 238.640 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 13.800 13.515 485.760 486.965 ;
      LAYER met1 ;
        RECT 0.070 13.360 493.050 487.120 ;
      LAYER met2 ;
        RECT 0.100 495.720 19.130 496.810 ;
        RECT 19.970 495.720 44.890 496.810 ;
        RECT 45.730 495.720 70.650 496.810 ;
        RECT 71.490 495.720 96.410 496.810 ;
        RECT 97.250 495.720 122.170 496.810 ;
        RECT 123.010 495.720 147.930 496.810 ;
        RECT 148.770 495.720 173.690 496.810 ;
        RECT 174.530 495.720 202.670 496.810 ;
        RECT 203.510 495.720 228.430 496.810 ;
        RECT 229.270 495.720 254.190 496.810 ;
        RECT 255.030 495.720 279.950 496.810 ;
        RECT 280.790 495.720 305.710 496.810 ;
        RECT 306.550 495.720 331.470 496.810 ;
        RECT 332.310 495.720 357.230 496.810 ;
        RECT 358.070 495.720 382.990 496.810 ;
        RECT 383.830 495.720 408.750 496.810 ;
        RECT 409.590 495.720 434.510 496.810 ;
        RECT 435.350 495.720 460.270 496.810 ;
        RECT 461.110 495.720 486.030 496.810 ;
        RECT 486.870 495.720 493.020 496.810 ;
        RECT 0.100 4.280 493.020 495.720 ;
        RECT 0.650 4.000 25.570 4.280 ;
        RECT 26.410 4.000 51.330 4.280 ;
        RECT 52.170 4.000 77.090 4.280 ;
        RECT 77.930 4.000 102.850 4.280 ;
        RECT 103.690 4.000 128.610 4.280 ;
        RECT 129.450 4.000 154.370 4.280 ;
        RECT 155.210 4.000 180.130 4.280 ;
        RECT 180.970 4.000 205.890 4.280 ;
        RECT 206.730 4.000 231.650 4.280 ;
        RECT 232.490 4.000 257.410 4.280 ;
        RECT 258.250 4.000 283.170 4.280 ;
        RECT 284.010 4.000 308.930 4.280 ;
        RECT 309.770 4.000 337.910 4.280 ;
        RECT 338.750 4.000 363.670 4.280 ;
        RECT 364.510 4.000 389.430 4.280 ;
        RECT 390.270 4.000 415.190 4.280 ;
        RECT 416.030 4.000 440.950 4.280 ;
        RECT 441.790 4.000 466.710 4.280 ;
        RECT 467.550 4.000 492.470 4.280 ;
      LAYER met3 ;
        RECT 4.400 492.640 496.000 493.505 ;
        RECT 4.000 483.840 496.000 492.640 ;
        RECT 4.000 482.440 495.600 483.840 ;
        RECT 4.000 466.840 496.000 482.440 ;
        RECT 4.400 465.440 496.000 466.840 ;
        RECT 4.000 456.640 496.000 465.440 ;
        RECT 4.000 455.240 495.600 456.640 ;
        RECT 4.000 439.640 496.000 455.240 ;
        RECT 4.400 438.240 496.000 439.640 ;
        RECT 4.000 429.440 496.000 438.240 ;
        RECT 4.000 428.040 495.600 429.440 ;
        RECT 4.000 412.440 496.000 428.040 ;
        RECT 4.400 411.040 496.000 412.440 ;
        RECT 4.000 402.240 496.000 411.040 ;
        RECT 4.000 400.840 495.600 402.240 ;
        RECT 4.000 385.240 496.000 400.840 ;
        RECT 4.400 383.840 496.000 385.240 ;
        RECT 4.000 375.040 496.000 383.840 ;
        RECT 4.000 373.640 495.600 375.040 ;
        RECT 4.000 358.040 496.000 373.640 ;
        RECT 4.400 356.640 496.000 358.040 ;
        RECT 4.000 347.840 496.000 356.640 ;
        RECT 4.000 346.440 495.600 347.840 ;
        RECT 4.000 327.440 496.000 346.440 ;
        RECT 4.400 326.040 496.000 327.440 ;
        RECT 4.000 320.640 496.000 326.040 ;
        RECT 4.000 319.240 495.600 320.640 ;
        RECT 4.000 300.240 496.000 319.240 ;
        RECT 4.400 298.840 496.000 300.240 ;
        RECT 4.000 293.440 496.000 298.840 ;
        RECT 4.000 292.040 495.600 293.440 ;
        RECT 4.000 273.040 496.000 292.040 ;
        RECT 4.400 271.640 496.000 273.040 ;
        RECT 4.000 266.240 496.000 271.640 ;
        RECT 4.000 264.840 495.600 266.240 ;
        RECT 4.000 245.840 496.000 264.840 ;
        RECT 4.400 244.440 496.000 245.840 ;
        RECT 4.000 239.040 496.000 244.440 ;
        RECT 4.000 237.640 495.600 239.040 ;
        RECT 4.000 218.640 496.000 237.640 ;
        RECT 4.400 217.240 496.000 218.640 ;
        RECT 4.000 211.840 496.000 217.240 ;
        RECT 4.000 210.440 495.600 211.840 ;
        RECT 4.000 191.440 496.000 210.440 ;
        RECT 4.400 190.040 496.000 191.440 ;
        RECT 4.000 184.640 496.000 190.040 ;
        RECT 4.000 183.240 495.600 184.640 ;
        RECT 4.000 164.240 496.000 183.240 ;
        RECT 4.400 162.840 496.000 164.240 ;
        RECT 4.000 157.440 496.000 162.840 ;
        RECT 4.000 156.040 495.600 157.440 ;
        RECT 4.000 137.040 496.000 156.040 ;
        RECT 4.400 135.640 496.000 137.040 ;
        RECT 4.000 126.840 496.000 135.640 ;
        RECT 4.000 125.440 495.600 126.840 ;
        RECT 4.000 109.840 496.000 125.440 ;
        RECT 4.400 108.440 496.000 109.840 ;
        RECT 4.000 99.640 496.000 108.440 ;
        RECT 4.000 98.240 495.600 99.640 ;
        RECT 4.000 82.640 496.000 98.240 ;
        RECT 4.400 81.240 496.000 82.640 ;
        RECT 4.000 72.440 496.000 81.240 ;
        RECT 4.000 71.040 495.600 72.440 ;
        RECT 4.000 55.440 496.000 71.040 ;
        RECT 4.400 54.040 496.000 55.440 ;
        RECT 4.000 45.240 496.000 54.040 ;
        RECT 4.000 43.840 495.600 45.240 ;
        RECT 4.000 28.240 496.000 43.840 ;
        RECT 4.400 26.840 496.000 28.240 ;
        RECT 4.000 18.040 496.000 26.840 ;
        RECT 4.000 16.640 495.600 18.040 ;
        RECT 4.000 13.435 496.000 16.640 ;
      LAYER met4 ;
        RECT 129.095 15.135 208.920 484.665 ;
        RECT 211.320 15.135 212.220 484.665 ;
        RECT 214.620 15.135 388.920 484.665 ;
        RECT 391.320 15.135 392.220 484.665 ;
        RECT 394.620 15.135 478.105 484.665 ;
  END
END mem
END LIBRARY

