// This is the unpowered netlist.
module core (clk,
    o_mem_write_M,
    rst,
    i_instr_ID,
    i_read_data_M,
    o_data_addr_M,
    o_funct3_MEM,
    o_pc_IF,
    o_write_data_M);
 input clk;
 output o_mem_write_M;
 input rst;
 input [31:0] i_instr_ID;
 input [31:0] i_read_data_M;
 output [31:0] o_data_addr_M;
 output [2:0] o_funct3_MEM;
 output [31:0] o_pc_IF;
 output [31:0] o_write_data_M;

 wire net485;
 wire net486;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ;
 wire \U_CONTROL_UNIT.i_branch_EX ;
 wire \U_CONTROL_UNIT.i_jump_EX ;
 wire \U_DATAPATH.U_EX_MEM.i_funct3_EX[0] ;
 wire \U_DATAPATH.U_EX_MEM.i_funct3_EX[1] ;
 wire \U_DATAPATH.U_EX_MEM.i_funct3_EX[2] ;
 wire \U_DATAPATH.U_EX_MEM.i_mem_write_EX ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[10] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[11] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[12] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[13] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[14] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[15] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[16] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[17] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[18] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[19] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[20] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[21] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[22] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[23] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[24] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[25] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[26] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[27] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[28] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[29] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[2] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[30] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[31] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[3] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[4] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[5] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[6] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[7] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[8] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[9] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[0] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[1] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[2] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[3] ;
 wire \U_DATAPATH.U_EX_MEM.i_reg_write_EX ;
 wire \U_DATAPATH.U_EX_MEM.i_result_src_EX[0] ;
 wire \U_DATAPATH.U_EX_MEM.i_result_src_EX[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[10] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[11] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[12] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[13] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[14] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[15] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[16] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[17] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[18] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[19] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[20] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[21] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[22] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[23] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[24] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[25] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[26] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[27] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[28] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[29] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[30] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[31] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[4] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[5] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[6] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[7] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[8] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[9] ;
 wire \U_DATAPATH.U_EX_MEM.o_mem_write_M ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[10] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[11] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[12] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[13] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[14] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[15] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[16] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[17] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[18] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[19] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[20] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[21] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[22] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[23] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[24] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[25] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[26] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[27] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[28] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[29] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[30] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[31] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[4] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[5] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[6] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[7] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[8] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[9] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[10] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[11] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[12] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[13] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[14] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[15] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[16] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[17] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[18] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[19] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[20] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[21] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[22] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[23] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[24] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[25] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[26] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[27] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[28] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[29] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[30] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[31] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[4] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[5] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[6] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[7] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[8] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[9] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_reg_write_M ;
 wire \U_DATAPATH.U_EX_MEM.o_result_src_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_result_src_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[10] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[11] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[12] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[13] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[14] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[15] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[16] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[17] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[18] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[19] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[20] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[21] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[22] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[23] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[24] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[25] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[26] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[27] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[28] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[29] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[30] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[31] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[4] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[5] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[6] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[7] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[8] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[9] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[0] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[1] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[0] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[1] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[0] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[1] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.o_addr_src_EX ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_src_EX ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[9] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[9] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[9] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[10] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[11] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[12] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[13] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[14] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[15] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[16] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[17] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[18] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[19] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[20] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[21] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[22] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[23] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[24] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[25] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[26] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[27] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[28] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[29] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[2] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[30] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[31] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[3] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[4] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[5] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[6] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[7] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[8] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[9] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[11] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[19] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[24] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[25] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[26] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[27] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[28] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[29] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[1] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[1] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[1] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net21;
 wire net210;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net211;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net212;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net213;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net216;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net217;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net218;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net219;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net22;
 wire net220;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net221;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net222;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net223;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net235;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net236;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net237;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net238;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net239;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net24;
 wire net240;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net2172));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net2240));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net2240));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net2240));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net2240));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net2240));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net2240));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net2283));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net2138));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__B (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__B (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__S0 (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__S1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A1 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__B1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__B (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__B1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A_N (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A_N (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__B1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__B2 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__A1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__B1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__B (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__B (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A_N (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__B1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A_N (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__B1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__B2 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__B (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__B (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__B (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A2 (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A2 (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__B (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__B (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__B1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__B1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__B1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__C (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A1 (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__B1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__B (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__B (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A1 (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__B1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A1 (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__C (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__B1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__B (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__B (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__A (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__B (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A_N (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__B1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__A1 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__B (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__B (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A_N (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__C (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__B (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__B (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__B (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__A1 (.DIODE(_1583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__B1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__B2 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A2 (.DIODE(net2141));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__B1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__B (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__B (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A_N (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__B1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__B2 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__B (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__A_N (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__B1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__B2 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A2 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__B1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__B (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__B (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A_N (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__C (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__B1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A1 (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__B (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__B (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A_N (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__B1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__B2 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A2 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__B1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__B (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__B (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A_N (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__B1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__B2 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__B1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__A (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__B (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__B (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__C (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__A1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__A2 (.DIODE(_1657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A2 (.DIODE(_1657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__B1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__B (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__B (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A1 (.DIODE(_1666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__C (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__B (.DIODE(net2333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__A1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__A2 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A2 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__B1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__B (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__B (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__A2 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__C (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__C (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A3 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__B1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__B1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__A2 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__C (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A0 (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A1 (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__B1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__A (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__B (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__B (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A_N (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__A1 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__B1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__A0 (.DIODE(net2184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__A1 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__B (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__A1 (.DIODE(_1715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__B (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__A1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__A2 (.DIODE(_1718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A2 (.DIODE(_1718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__B (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__C (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__B (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__B (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__B (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__B (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__B (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__B (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__B (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__B (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__C (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__B (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__C (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__B1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__B1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__C (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__A1 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__B1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A_N (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__B (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__C (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__A1 (.DIODE(_1759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__B1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__B (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__B (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__B1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A1 (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__B (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__B (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__A_N (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__A1 (.DIODE(_1776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__B1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__B2 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A2 (.DIODE(_1779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__B (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__A_N (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__C (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__B1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__A1 (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__C (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__B (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__B (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__A_N (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4149__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__C (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__A1 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__B1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__B (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__C (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__B1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A1 (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__A2 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__B (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__B (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__A1 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__B2 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__A1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__A2 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__B (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__C (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__B (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__A_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__A1 (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__B (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__C (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__B2 (.DIODE(_1464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__A (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__B (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__A (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__B (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__A (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A_N (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__A_N (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__C1 (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__A_N (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__B1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__B (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__A (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__A_N (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__A_N (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__B (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__A_N (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__A_N (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__A3 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__B1 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__A_N (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__B (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__B1 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__A2 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__B1 (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__A_N (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__B (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__A_N (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__B (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__A2 (.DIODE(_1881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__A_N (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__A_N (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__B (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4237__A_N (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__A_N (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__A3 (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__B1 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__A_N (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__B (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__A2 (.DIODE(_1875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__A3 (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__A (.DIODE(net2333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__B (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__C (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__A (.DIODE(net2333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__B (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__S (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A_N (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__B (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__B1_N (.DIODE(_1938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__C_N (.DIODE(_1938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__A_N (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__S (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A2 (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__B (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__A (.DIODE(_1943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__A (.DIODE(net2184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__S (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__S (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__S (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__S (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__S (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__S (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__A0 (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__S (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__A (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__S (.DIODE(net2257));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__A1 (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__B (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__S (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__B1_N (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__C_N (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A_N (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__B (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__C (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__S (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__A2 (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__B (.DIODE(_2085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__S (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__A (.DIODE(_2090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__S (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__B (.DIODE(_2100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__B (.DIODE(_2100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__S (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__S (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__S (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__B (.DIODE(_2108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__S (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__S (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__S (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__S (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__S (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__B (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__S (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__S (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__A1 (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__S (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__A (.DIODE(_2153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__S (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__S (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__A (.DIODE(_2153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__S (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__S (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__S (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__A (.DIODE(_2180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__S (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__A (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__A (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__B (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__B (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__A (.DIODE(_2178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A (.DIODE(_2178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A1 (.DIODE(_2178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__B1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A (.DIODE(_2153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A (.DIODE(_2153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A1 (.DIODE(_2090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A3 (.DIODE(_2108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__B (.DIODE(_2108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__A2 (.DIODE(_2108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__B1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A (.DIODE(_2090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__A1 (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__A3 (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__B1 (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__A (.DIODE(_2090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__A (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__B (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__S (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A1 (.DIODE(net2014));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__A (.DIODE(_1943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A1 (.DIODE(net2014));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__B (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__B (.DIODE(\U_DATAPATH.U_EX_MEM.o_write_data_M[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__S (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__S (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__S (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__S (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__S (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__A1 (.DIODE(_2108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__S (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A0 (.DIODE(net2080));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A1 (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__S (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A1 (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__S (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__S (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__A0 (.DIODE(net2041));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__S (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__A0 (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__S (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__S (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__A1 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__S1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__S0 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__S1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__S0 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__S1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__S1 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__S0 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__S1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__S0 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__S1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__S1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__S1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__S1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__S1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__S0 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__S1 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__S1 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__S0 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__S1 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__S0 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__S1 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__S0 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__S0 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__S0 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__S1 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__S0 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__S0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__S0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__S1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__S1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__S0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__S1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__S0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__S1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__S1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__S1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__S0 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__S1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__S0 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__S1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__S1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__S0 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__S0 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__S1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__S1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__S1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__S1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__S1 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__S1 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__S1 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__S1 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__S0 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__S0 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__S1 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__S0 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__S1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__S1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__S1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__S0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__S1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__S0 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__S0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__S1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__S (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__C_N (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__B (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__B (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A (.DIODE(net2086));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A1 (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__B (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__S (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__C_N (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__S (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__C_N (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A (.DIODE(net2128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A (.DIODE(net2103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A (.DIODE(net2134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__A (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A (.DIODE(net2055));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A (.DIODE(net2105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A (.DIODE(net2172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__B (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A (.DIODE(net1997));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A (.DIODE(net2214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A (.DIODE(net2007));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A (.DIODE(net2138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A (.DIODE(net2190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A (.DIODE(net2019));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__B (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A1 (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A1 (.DIODE(net2041));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A1 (.DIODE(net2080));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__C1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__A1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__A1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__A1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A2 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__A2 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A (.DIODE(net2055));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__B (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__C (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A_N (.DIODE(net2055));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__B (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__B (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__B (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A (.DIODE(net2055));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A (.DIODE(net2055));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__B (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__B (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__C_N (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A1 (.DIODE(net2055));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A2 (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__B (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A1 (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A2 (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A (.DIODE(net2240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__C (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A (.DIODE(net2055));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__C (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__C (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__C (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__C (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A (.DIODE(net2086));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__B (.DIODE(net2044));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__C (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__C (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__C (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__C (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__C (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__C (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__C (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__B (.DIODE(net2044));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__C (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__C (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__C (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__C (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__B (.DIODE(net2044));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__C (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__C (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__C (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__C (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__C (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__C (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__C (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__C (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__C (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__C (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__C (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__C (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__C (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__C (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__C (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__C (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A (.DIODE(net2128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A (.DIODE(net2103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A (.DIODE(net2134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A2 (.DIODE(net2257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__B (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__B (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__B (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A0 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A1 (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A2 (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A0 (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A1 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A2 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A3 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__S0 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A0 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A1 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A0 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A1 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A2 (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A3 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__A0 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__A1 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__A0 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__A1 (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A0 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A1 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A0 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A1 (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A0 (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A1 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A0 (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A1 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A1 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A0 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A1 (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__A1 (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__B (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__B (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__C (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__D (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__B1 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__B (.DIODE(_2864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__B (.DIODE(_2864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__C (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__C1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__B2 (.DIODE(_2853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__C1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A0 (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A1 (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A2 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A3 (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__A1 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A1 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A2 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A3 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A0 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A2 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A3 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A0 (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5913__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A1 (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A1 (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A1 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__B2 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__C (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__B1 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A0 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A1 (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__B2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__C1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A1 (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A1_N (.DIODE(_2853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__B2 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A0 (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A2 (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A3 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A0 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A2 (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A3 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A0 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A1 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A0 (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A0 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A0 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A2 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A3 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__B (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__A0 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A0 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A1 (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A2 (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A3 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__S0 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A0 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A1 (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A2 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A3 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__S0 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__A2 (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__B (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__A (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__B1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__A2 (.DIODE(_2857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__B1 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__C1 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__A2 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__C1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__C1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A0 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A1 (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A2 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A3 (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A0 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A1 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A2 (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A3 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__A0 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__A1 (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__A2 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__A (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__S (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__S (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__A1 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__B2 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__A (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__B (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__A (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__A (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__A (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__A0 (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__A1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__A (.DIODE(_2853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__C1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A1 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A0 (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A1 (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A2 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A3 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A0 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A1 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A2 (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A3 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__S (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__S (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__A2 (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__B (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6026__A (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__A (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__A1 (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__S (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__A2 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A0 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A1 (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A3 (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__C1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__A1 (.DIODE(_2853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__C1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__C1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__A (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__C1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__A0 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__A1 (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A1 (.DIODE(_2864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__B1 (.DIODE(_3027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__C1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__A (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__B1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A2 (.DIODE(_2857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__B1 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__C1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A0 (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A1 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A2 (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A3 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__B (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__C1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__A (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A0 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A1 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A2 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A3 (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__A2 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__B1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A1_N (.DIODE(_2864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__A1 (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__A (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__C1 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__C1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__A (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__A (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A0 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A1 (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A2 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A3 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__B2 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__C1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A2 (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__A (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A0 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A1 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A2 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A3 (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__A2 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__C1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A2 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__C1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__A (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A0 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A1 (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A2 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A3 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__C1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__A2 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__C1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__A (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__A (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__B1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A0 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A1 (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A2 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A3 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__C1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__B2 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__C1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6228__A (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A1 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__B1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__A1 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__A0 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__A2 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__A3 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6237__C1 (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A1_N (.DIODE(_2864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__B2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__B2 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__A2 (.DIODE(_3199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__D1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__C1 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__A (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__A (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__A1 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A0 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A1 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A2 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A3 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__A2 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__B1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__A1 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__B2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__A1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__B1 (.DIODE(_3218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__A2 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__C1 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__A (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__A (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A0 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A2 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A3 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__A1_N (.DIODE(_2864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__B2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__B2 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__A2 (.DIODE(_3235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__C1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__A1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__B1 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__C1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__A (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__A (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__A (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A0 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A2 (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A3 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__B2 (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__C1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A1 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__B1 (.DIODE(_3253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__A1 (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__B1 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A1 (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__B1 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__S (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A1 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__B1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__A3 (.DIODE(_3261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__B (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__A1 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__A2 (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__A3 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__C1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__B1 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A2 (.DIODE(_3276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__D1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__C1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A2 (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A3 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__C1 (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__C1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__A2 (.DIODE(_3276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__B2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__B2 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__C1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__A (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__A (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__A (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__B1 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__C1 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__A2 (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__B1 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__B2 (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__C1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__A1 (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__A2 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A1 (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__A1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__B2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__B1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__A (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__A (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__A1 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__A3 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__S0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__C1 (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__B2 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__C1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A2 (.DIODE(_3276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__B2 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__A1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__B2 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A1 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__C1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__A (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__A (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A (.DIODE(_3333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A0 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A1 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A2 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__B1 (.DIODE(_3276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__B1 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__C1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__A2 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__C1 (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__A1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__C1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__A (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__A (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__A (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A1 (.DIODE(_3333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__A2 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__C1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__B2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__A0 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__A1 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__A2 (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__A3 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__A1_N (.DIODE(_2853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__B1 (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__A2 (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__C1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__A (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__A (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__A (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__A0 (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__A1 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__A2 (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__A3 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A1 (.DIODE(_2853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__C1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__C1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__B1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__B1 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__A2 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__C1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__A (.DIODE(_2864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A0 (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A1 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A2 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A3 (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__A1 (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__B1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__C1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__A (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__A (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6461__A (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A0 (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A1 (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A2 (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A3 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__S0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__A1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__B1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__A2 (.DIODE(_2864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__A (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__A (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__B1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A0 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A1 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A2 (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A3 (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__S0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__A1_N (.DIODE(_2853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A2 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__C1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__A1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__A2 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__C1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6498__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__A (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__A1 (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__A2 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__A3 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__A1_N (.DIODE(_2853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__A1_N (.DIODE(_2864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__B2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__C1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__A1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__C1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__A (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__A (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__A (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A0 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A1 (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A2 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A3 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__B2 (.DIODE(_2853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__B1 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__A1 (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__B1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__A1 (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__A2 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A1 (.DIODE(_2864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__A1 (.DIODE(_1647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__A2 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__C1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__A (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__A (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__A0 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__A1 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__A2 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__A3 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__B1 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__C1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6544__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__A3 (.DIODE(_3276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6547__A2 (.DIODE(_3480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6547__C1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__A (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__A (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__A0 (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__A1 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__A2 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__A3 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__B2 (.DIODE(_2853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__A2 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__C1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__A1 (.DIODE(_2864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__B1 (.DIODE(_3495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__A2 (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__B (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A0 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A2 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A3 (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__S0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__B2 (.DIODE(_2853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__B1 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__C1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__C1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A0 (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A2 (.DIODE(_1503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A3 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A2 (.DIODE(_3253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__C1 (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A2 (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__B1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__A1 (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__A2 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__C1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__A3 (.DIODE(_3276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__A2 (.DIODE(_1467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__C1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__B (.DIODE(_1697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A3 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__B1 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__B (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__B (.DIODE(_1718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__B1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__B (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__B (.DIODE(_1779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__B (.DIODE(_1759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__B (.DIODE(net2174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__B (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__B (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__B (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__B (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__B (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__B (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__B1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__B (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__B (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__B (.DIODE(net2141));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__B (.DIODE(net2304));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__B (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__B (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__B (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__B (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__B (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__B (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__B (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__A (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__C (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__A (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__A (.DIODE(net2055));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__C (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__A1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__A1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__A2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__C (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A3 (.DIODE(_3540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__B (.DIODE(_3540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__A3 (.DIODE(_3540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__A1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__A1 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__A1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__A1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__6842__A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__6845__A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__6845__B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6846__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6862__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6862__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__A1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__B1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__A1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__A1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__A1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6924__A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__6924__C (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6926__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__A1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__B (.DIODE(_3583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__A3 (.DIODE(_3583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__A1 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__A1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__A1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__A1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6948__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6958__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6958__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6962__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6962__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6964__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6964__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__A1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__A3 (.DIODE(_3583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6968__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6968__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6976__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6976__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6978__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__6978__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6981__A3 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6984__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__6984__B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6988__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6990__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6990__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6992__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6992__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6998__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6998__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__A1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__7009__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__7009__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7009__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7012__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__7012__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7012__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7016__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__7016__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7016__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7017__A1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__7017__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7017__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7020__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__7020__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7022__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__7022__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7022__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7023__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__7024__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7029__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7029__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7033__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__7033__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7033__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__A1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7041__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__7041__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7041__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7048__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__7048__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7048__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__A1 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7058__A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__7058__C (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7059__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__7059__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7060__A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__7060__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7061__A1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7061__A3 (.DIODE(_3625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__A1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7065__A1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7065__A3 (.DIODE(_3625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__A1 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7072__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__7072__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7074__A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__7074__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__A1 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__A1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7082__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__7082__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7085__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__7085__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__A1 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7093__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7093__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7098__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__7098__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7102__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__7102__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7105__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__7105__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7109__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__7109__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__A1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__A3 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__A1 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7118__A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__7118__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7119__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__7119__A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__C (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__A (.DIODE(_1679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__A (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__A1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__A3 (.DIODE(_3659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7128__A (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7128__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7129__A1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7129__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7130__A (.DIODE(_1716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7130__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__A1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7133__A2 (.DIODE(_3659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7136__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7137__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__7137__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7139__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__7139__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7140__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__A1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7146__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7147__A1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7147__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7148__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__7148__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7149__A1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__7149__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7150__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7152__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7153__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7153__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7155__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__7155__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7159__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7159__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7161__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__7161__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7164__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__7164__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7165__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__7165__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7166__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7168__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__7168__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7170__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7171__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__7171__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7173__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__7173__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7174__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__7174__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__A1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7179__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__7179__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7183__A1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__7183__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7185__A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7186__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7187__A (.DIODE(net2055));
 sky130_fd_sc_hd__diode_2 ANTENNA__7187__B (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__7187__C (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA__7189__A1_N (.DIODE(net2190));
 sky130_fd_sc_hd__diode_2 ANTENNA__7192__A1 (.DIODE(net2190));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__A1 (.DIODE(net2190));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__A2 (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__C1 (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__7198__A1 (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7198__B2 (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7202__A1 (.DIODE(net2190));
 sky130_fd_sc_hd__diode_2 ANTENNA__7204__A0 (.DIODE(net2190));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__A (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__A1 (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__B2 (.DIODE(net2206));
 sky130_fd_sc_hd__diode_2 ANTENNA__7211__A0 (.DIODE(net2190));
 sky130_fd_sc_hd__diode_2 ANTENNA__7212__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7213__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7214__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__7215__A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__7216__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7217__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7218__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7219__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__7220__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__7223__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__7225__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__7227__A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__7229__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__7230__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__7231__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__7232__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__7233__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__7234__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__7235__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__7236__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__7239__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__7240__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__7241__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__7242__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__7243__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__7245__A (.DIODE(net2019));
 sky130_fd_sc_hd__diode_2 ANTENNA__7245__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__7245__C (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__7246__A (.DIODE(net2019));
 sky130_fd_sc_hd__diode_2 ANTENNA__7247__A (.DIODE(net2190));
 sky130_fd_sc_hd__diode_2 ANTENNA__7247__B (.DIODE(net2074));
 sky130_fd_sc_hd__diode_2 ANTENNA__7248__A1 (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA__7248__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7249__A (.DIODE(net2138));
 sky130_fd_sc_hd__diode_2 ANTENNA__7249__B (.DIODE(net2074));
 sky130_fd_sc_hd__diode_2 ANTENNA__7250__A1 (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA__7250__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7251__A (.DIODE(net2007));
 sky130_fd_sc_hd__diode_2 ANTENNA__7251__B (.DIODE(net2074));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__A1 (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__A (.DIODE(net2214));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__B (.DIODE(net2074));
 sky130_fd_sc_hd__diode_2 ANTENNA__7254__A1 (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA__7254__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__A (.DIODE(net1997));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__B (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7256__A1 (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA__7256__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__B (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7258__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7259__A (.DIODE(net2172));
 sky130_fd_sc_hd__diode_2 ANTENNA__7259__B (.DIODE(net2074));
 sky130_fd_sc_hd__diode_2 ANTENNA__7260__A1 (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA__7260__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7261__A (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__7261__B (.DIODE(net2074));
 sky130_fd_sc_hd__diode_2 ANTENNA__7262__A1 (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA__7262__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7263__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__7263__B (.DIODE(net2074));
 sky130_fd_sc_hd__diode_2 ANTENNA__7264__A1 (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA__7264__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7265__A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__7265__B (.DIODE(net2074));
 sky130_fd_sc_hd__diode_2 ANTENNA__7266__A1 (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA__7266__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7267__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__7267__B (.DIODE(net2074));
 sky130_fd_sc_hd__diode_2 ANTENNA__7268__A1 (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA__7268__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7269__A (.DIODE(net2105));
 sky130_fd_sc_hd__diode_2 ANTENNA__7269__B (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7270__A (.DIODE(net2019));
 sky130_fd_sc_hd__diode_2 ANTENNA__7271__A2 (.DIODE(_3727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7271__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7272__A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__7272__B (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7273__A1 (.DIODE(_3727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7273__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7274__A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__7274__B (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7275__A1 (.DIODE(_3727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7275__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7276__A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__7276__B (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7277__A1 (.DIODE(_3727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7277__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7278__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__7278__B (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7279__A1 (.DIODE(_3727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7279__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7280__A (.DIODE(net2055));
 sky130_fd_sc_hd__diode_2 ANTENNA__7280__B (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7281__A1 (.DIODE(_3727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7281__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7282__A (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__7282__B (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7283__A1 (.DIODE(_3727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7283__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7284__A (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA__7284__B (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7285__A1 (.DIODE(_3727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7285__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7286__B (.DIODE(_3727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7287__A1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__7287__B2 (.DIODE(net2128));
 sky130_fd_sc_hd__diode_2 ANTENNA__7289__A (.DIODE(net2190));
 sky130_fd_sc_hd__diode_2 ANTENNA__7290__A (.DIODE(net2138));
 sky130_fd_sc_hd__diode_2 ANTENNA__7291__A (.DIODE(net2007));
 sky130_fd_sc_hd__diode_2 ANTENNA__7292__A (.DIODE(net2214));
 sky130_fd_sc_hd__diode_2 ANTENNA__7293__A (.DIODE(net1997));
 sky130_fd_sc_hd__diode_2 ANTENNA__7295__A (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7295__B (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7296__A1 (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7296__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7297__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7297__B1 (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7297__B2 (.DIODE(net2172));
 sky130_fd_sc_hd__diode_2 ANTENNA__7298__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__7298__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7299__A1 (.DIODE(net2134));
 sky130_fd_sc_hd__diode_2 ANTENNA__7299__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7299__B1 (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7299__B2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__7300__A (.DIODE(net2044));
 sky130_fd_sc_hd__diode_2 ANTENNA__7301__A1 (.DIODE(net2103));
 sky130_fd_sc_hd__diode_2 ANTENNA__7301__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7301__B1 (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7301__B2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__7302__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__7303__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7303__B1 (.DIODE(_3738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7303__B2 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__7304__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__7305__A1 (.DIODE(net2128));
 sky130_fd_sc_hd__diode_2 ANTENNA__7305__A3 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7305__B2 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__7306__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__7306__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7311__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__7312__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__7313__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__7314__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__7315__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__7316__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__7317__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__7318__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__7319__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__7320__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__7321__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__7322__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__7323__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__7324__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__7325__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__7326__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__7327__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__7328__A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__7329__A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__7330__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__7331__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__7332__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__7333__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__7334__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__7335__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__7336__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__7337__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__7338__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__7339__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__7356__18_A (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7358__20_A (.DIODE(clknet_leaf_33_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7360__22_A (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7367__29_A (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7379__41_A (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7382__44_A (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7391__53_A (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7392__54_A (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7396__58_A (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7397__59_A (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7399__61_A (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7401__63_A (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7403__65_A (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7404__66_A (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7405__67_A (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7414__76_A (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7416__78_A (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7421__83_A (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7428__90_A (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7431__93_A (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7432__94_A (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7434__96_A (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7435__97_A (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7452__114_A (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7453__115_A (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7455__117_A (.DIODE(clknet_leaf_33_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7456__118_A (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7464__126_A (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7468__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__7469__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__7470__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__7471__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__7472__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__7473__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__7474__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__7475__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__7476__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__7477__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__7478__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__7479__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__7480__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__7481__A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__7482__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__7483__A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__7484__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__7485__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__7486__A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__7487__A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__7488__A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__7489__A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__7490__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__7491__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__7492__A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__7493__A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__7494__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__7495__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__7496__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__7497__A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__7500__RESET_B (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7508__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7519__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7526__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7527__CLK (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7528__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7538__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7539__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7540__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7551__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7555__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7556__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7557__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7558__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7561__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7562__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7563__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7564__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7569__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7570__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7574__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7576__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7582__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7583__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7589__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7598__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7615__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7617__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7631__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7639__CLK (.DIODE(clknet_leaf_33_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7640__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7651__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7655__CLK (.DIODE(clknet_leaf_33_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7663__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7669__CLK (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7704__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7710__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7715__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7756__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7759__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7765__CLK (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7768__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7774__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7776__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7778__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7779__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7788__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7791__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7797__CLK (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7806__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7808__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7810__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7811__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7823__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7832__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7843__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7846__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7847__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7848__D (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7857__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7858__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7859__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7871__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7873__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7875__CLK (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7876__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7885__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7888__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7897__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7904__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7934__CLK (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7965__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7966__CLK (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7982__D (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7994__D (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7998__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7999__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8004__D (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8014__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8016__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8017__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8018__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8032__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8033__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8034__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8046__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8050__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8051__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8055__CLK (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8070__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8071__CLK (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8076__CLK (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8076__D (.DIODE(_0836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8078__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8081__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8085__CLK (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8086__D (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8089__D (.DIODE(_0849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8090__D (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8097__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8100__CLK (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8109__CLK (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8110__CLK (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8114__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8115__CLK (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8116__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8116__D (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8117__CLK (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8118__D (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8120__D (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8121__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8126__CLK (.DIODE(clknet_leaf_33_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8127__CLK (.DIODE(clknet_leaf_33_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8128__CLK (.DIODE(clknet_leaf_33_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8129__CLK (.DIODE(clknet_leaf_33_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8138__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8139__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8144__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8149__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8151__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8153__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8157__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8159__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8161__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8170__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8176__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8183__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8184__CLK (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8185__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8187__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8189__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8191__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8192__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8206__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8207__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8213__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8215__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8219__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8220__CLK (.DIODE(clknet_leaf_74_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8221__D (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8222__D (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8256__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8257__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8266__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8268__CLK (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8273__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8280__CLK (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8283__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8284__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8286__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8287__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8289__D (.DIODE(_1017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8291__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8359__CLK (.DIODE(clknet_leaf_33_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8366__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8372__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8373__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8382__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8397__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8399__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8404__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8416__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8418__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8426__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8431__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8448__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8459__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8463__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8469__CLK (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8478__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8510__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8515__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8519__CLK (.DIODE(clknet_leaf_33_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8527__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8533__CLK (.DIODE(clknet_leaf_47_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8542__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8547__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8551__CLK (.DIODE(clknet_leaf_33_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8556__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8565__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8574__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8579__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8588__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8589__CLK (.DIODE(clknet_leaf_3_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8602__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8605__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8606__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8607__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8608__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8613__CLK (.DIODE(clknet_leaf_33_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8620__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8621__CLK (.DIODE(clknet_leaf_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8627__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8641__CLK (.DIODE(clknet_leaf_54_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8651__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8652__CLK (.DIODE(clknet_leaf_4_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8658__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8688__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8692__CLK (.DIODE(clknet_leaf_42_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8695__CLK (.DIODE(clknet_leaf_52_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8698__CLK (.DIODE(clknet_leaf_33_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8707__CLK (.DIODE(clknet_leaf_71_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8715__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__8718__CLK (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(_1721_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(_1721_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(_3622_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(_3622_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(_3580_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(_3580_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(_3575_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(_3575_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(_2770_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(_2770_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(_2750_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(_2750_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(_3659_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(_3625_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(_3618_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(_3618_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(_3583_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(_3582_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(_3582_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(_2754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(_2754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_A (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_A (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(_1464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(_1464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(_3616_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout311_A (.DIODE(_3616_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout312_A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout313_A (.DIODE(_3540_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout316_A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout319_A (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(_1716_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout331_A (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout332_A (.DIODE(_1679_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout333_A (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout334_A (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout349_A (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout350_A (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout351_A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout353_A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout356_A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout358_A (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout359_A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout361_A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout362_A (.DIODE(_2857_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout363_A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout364_A (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout366_A (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout367_A (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout377_A (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout381_A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout382_A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout384_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout385_A (.DIODE(net2256));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout386_A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout387_A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout388_A (.DIODE(net2256));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout389_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout390_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout391_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout392_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout393_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout394_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout395_A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout396_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout397_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout399_A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout400_A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout401_A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout402_A (.DIODE(net2166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout403_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout404_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout405_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout406_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout407_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout408_A (.DIODE(net2166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout409_A (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout410_A (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout411_A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout412_A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout413_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout414_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout415_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout416_A (.DIODE(net2181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout417_A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout418_A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout419_A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout420_A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout421_A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout422_A (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout423_A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout424_A (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout425_A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout427_A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout428_A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout429_A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout430_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout431_A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout432_A (.DIODE(net2143));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout433_A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout434_A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout435_A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout436_A (.DIODE(net2143));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout437_A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout438_A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout439_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout440_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout441_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout442_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout443_A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout444_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout445_A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout446_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout447_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout448_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout449_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout450_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout451_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout452_A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout453_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout454_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout455_A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout456_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout457_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout458_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout459_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout460_A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout461_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout462_A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout463_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout464_A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout465_A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout466_A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout467_A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout468_A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout469_A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout470_A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout471_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout473_A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout474_A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout475_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout476_A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout477_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout478_A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout479_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout480_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout481_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1393_A (.DIODE(net2206));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1397_A (.DIODE(_1943_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1409_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1419_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1420_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1424_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1429_A (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1434_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1436_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1438_A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1446_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1447_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1451_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1452_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1454_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1457_A (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1458_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1459_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1460_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1461_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1463_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1464_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1465_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1466_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1471_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1472_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1473_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1478_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1479_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1480_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1482_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1487_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1488_A (.DIODE(\U_DATAPATH.U_IF_ID.o_instr_ID[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1494_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1499_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1500_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1504_A (.DIODE(_1657_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1526_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1533_A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1549_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1555_A (.DIODE(\U_DATAPATH.U_IF_ID.o_instr_ID[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1557_A (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1564_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1589_A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1597_A (.DIODE(net2406));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1598_A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1618_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1623_A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1635_A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1639_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1666_A (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1687_A (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1693_A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1703_A (.DIODE(_1783_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1704_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1706_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1714_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1719_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1730_A (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1732_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1733_A (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1740_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1741_A (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1744_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1745_A (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1747_A (.DIODE(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1750_A (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1788_A (.DIODE(\U_DATAPATH.U_IF_ID.o_instr_ID[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap303_A (.DIODE(_2205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_output152_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_split1_A (.DIODE(net184));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _3754_ (.A(net480),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _3755_ (.A(net2194),
    .Y(_1407_));
 sky130_fd_sc_hd__inv_2 _3756_ (.A(net2073),
    .Y(_1408_));
 sky130_fd_sc_hd__inv_2 _3757_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .Y(_1409_));
 sky130_fd_sc_hd__inv_2 _3758_ (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ),
    .Y(_1410_));
 sky130_fd_sc_hd__inv_2 _3759_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .Y(_1411_));
 sky130_fd_sc_hd__inv_2 _3760_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .Y(_1412_));
 sky130_fd_sc_hd__inv_2 _3761_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .Y(_1413_));
 sky130_fd_sc_hd__inv_2 _3762_ (.A(net380),
    .Y(_1414_));
 sky130_fd_sc_hd__inv_2 _3763_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .Y(_1415_));
 sky130_fd_sc_hd__inv_2 _3764_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ),
    .Y(_1416_));
 sky130_fd_sc_hd__inv_2 _3765_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ),
    .Y(_1417_));
 sky130_fd_sc_hd__inv_2 _3766_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ),
    .Y(_1418_));
 sky130_fd_sc_hd__inv_2 _3767_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ),
    .Y(_1419_));
 sky130_fd_sc_hd__inv_2 _3768_ (.A(net1507),
    .Y(_1420_));
 sky130_fd_sc_hd__inv_2 _3769__1 (.A(clknet_leaf_37_clk),
    .Y(net489));
 sky130_fd_sc_hd__nand2b_1 _3770_ (.A_N(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .Y(_1421_));
 sky130_fd_sc_hd__and2b_1 _3771_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .B(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .X(_1422_));
 sky130_fd_sc_hd__nand2b_1 _3772_ (.A_N(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .Y(_1423_));
 sky130_fd_sc_hd__nor4_1 _3773_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .C(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .D(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .Y(_1424_));
 sky130_fd_sc_hd__a221o_1 _3774_ (.A1(_1409_),
    .A2(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .B1(_1410_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .C1(_1422_),
    .X(_1425_));
 sky130_fd_sc_hd__nand2_1 _3775_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .Y(_1426_));
 sky130_fd_sc_hd__or2_1 _3776_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .X(_1427_));
 sky130_fd_sc_hd__a21o_1 _3777_ (.A1(_1426_),
    .A2(_1427_),
    .B1(_1424_),
    .X(_1428_));
 sky130_fd_sc_hd__o2111ai_2 _3778_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .A2(_1410_),
    .B1(_1421_),
    .C1(_1423_),
    .D1(net731),
    .Y(_1429_));
 sky130_fd_sc_hd__nor3_2 _3779_ (.A(_1425_),
    .B(_1428_),
    .C(_1429_),
    .Y(_1430_));
 sky130_fd_sc_hd__or3_1 _3780_ (.A(_1425_),
    .B(_1428_),
    .C(_1429_),
    .X(_1431_));
 sky130_fd_sc_hd__nand2b_1 _3781_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .Y(_1432_));
 sky130_fd_sc_hd__and2b_1 _3782_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .X(_1433_));
 sky130_fd_sc_hd__nand2b_1 _3783_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .Y(_1434_));
 sky130_fd_sc_hd__nand2_1 _3784_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .Y(_1435_));
 sky130_fd_sc_hd__or2_1 _3785_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .X(_1436_));
 sky130_fd_sc_hd__a21o_1 _3786_ (.A1(_1435_),
    .A2(_1436_),
    .B1(_1424_),
    .X(_1437_));
 sky130_fd_sc_hd__a221o_1 _3787_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .A2(_1411_),
    .B1(_1413_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .C1(_1433_),
    .X(_1438_));
 sky130_fd_sc_hd__o2111a_1 _3788_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .A2(_1411_),
    .B1(_1432_),
    .C1(_1434_),
    .D1(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .X(_1439_));
 sky130_fd_sc_hd__nor3b_2 _3789_ (.A(_1437_),
    .B(_1438_),
    .C_N(_1439_),
    .Y(_1440_));
 sky130_fd_sc_hd__or3b_4 _3790_ (.A(_1437_),
    .B(_1438_),
    .C_N(_1439_),
    .X(_1441_));
 sky130_fd_sc_hd__nor2_8 _3791_ (.A(net355),
    .B(_1441_),
    .Y(_1442_));
 sky130_fd_sc_hd__nor2_8 _3792_ (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(net438),
    .Y(_1443_));
 sky130_fd_sc_hd__or2_2 _3793_ (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(net437),
    .X(_1444_));
 sky130_fd_sc_hd__and2_2 _3794_ (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(net437),
    .X(_1445_));
 sky130_fd_sc_hd__mux4_2 _3795_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[31] ),
    .A1(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[31] ),
    .A2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[31] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[31] ),
    .S0(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .S1(net437),
    .X(_1446_));
 sky130_fd_sc_hd__nor2_2 _3796_ (.A(net356),
    .B(net351),
    .Y(_1447_));
 sky130_fd_sc_hd__a22o_1 _3797_ (.A1(_1442_),
    .A2(_1446_),
    .B1(net308),
    .B2(net2003),
    .X(_1448_));
 sky130_fd_sc_hd__a21oi_2 _3798_ (.A1(net623),
    .A2(net356),
    .B1(net2004),
    .Y(_1449_));
 sky130_fd_sc_hd__nand2_1 _3799_ (.A(net2269),
    .B(net379),
    .Y(_1450_));
 sky130_fd_sc_hd__o21ai_4 _3800_ (.A1(net379),
    .A2(_1449_),
    .B1(_1450_),
    .Y(_1451_));
 sky130_fd_sc_hd__or4_1 _3801_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ),
    .C(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ),
    .D(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ),
    .X(_1452_));
 sky130_fd_sc_hd__o2bb2a_4 _3802_ (.A1_N(_1418_),
    .A2_N(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .B1(_1410_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .X(_1453_));
 sky130_fd_sc_hd__o22a_1 _3803_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .A2(_1417_),
    .B1(_1418_),
    .B2(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .X(_1454_));
 sky130_fd_sc_hd__a22oi_1 _3804_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .A2(_1416_),
    .B1(_1417_),
    .B2(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .Y(_1455_));
 sky130_fd_sc_hd__o211a_1 _3805_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .A2(_1416_),
    .B1(_1452_),
    .C1(\U_DATAPATH.U_EX_MEM.o_reg_write_M ),
    .X(_1456_));
 sky130_fd_sc_hd__o2111a_4 _3806_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ),
    .A2(_1415_),
    .B1(_1454_),
    .C1(_1455_),
    .D1(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__and2b_1 _3807_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .X(_1458_));
 sky130_fd_sc_hd__a221o_1 _3808_ (.A1(_1411_),
    .A2(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ),
    .B1(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ),
    .B2(_1413_),
    .C1(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__xor2_1 _3809_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ),
    .X(_1460_));
 sky130_fd_sc_hd__a221o_1 _3810_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .A2(_1416_),
    .B1(_1418_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .C1(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__o211a_1 _3811_ (.A1(_1412_),
    .A2(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .B1(_1452_),
    .C1(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .X(_1462_));
 sky130_fd_sc_hd__or3b_2 _3812_ (.A(_1459_),
    .B(_1461_),
    .C_N(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__a21oi_4 _3813_ (.A1(net366),
    .A2(net349),
    .B1(_1463_),
    .Y(_1464_));
 sky130_fd_sc_hd__and3_1 _3814_ (.A(net623),
    .B(net367),
    .C(net350),
    .X(_1465_));
 sky130_fd_sc_hd__a21boi_4 _3815_ (.A1(net366),
    .A2(net349),
    .B1_N(_1463_),
    .Y(_1466_));
 sky130_fd_sc_hd__a221o_4 _3816_ (.A1(net370),
    .A2(net307),
    .B1(net305),
    .B2(net2351),
    .C1(_1465_),
    .X(_1467_));
 sky130_fd_sc_hd__inv_2 _3817_ (.A(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__xnor2_2 _3818_ (.A(_1451_),
    .B(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__and2b_1 _3819_ (.A_N(net437),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[28] ),
    .X(_1470_));
 sky130_fd_sc_hd__and2b_1 _3820_ (.A_N(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(net437),
    .X(_1471_));
 sky130_fd_sc_hd__a221o_1 _3821_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[28] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[28] ),
    .C1(_1470_),
    .X(_1472_));
 sky130_fd_sc_hd__mux2_1 _3822_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[28] ),
    .A1(_1472_),
    .S(net373),
    .X(_1473_));
 sky130_fd_sc_hd__a22o_1 _3823_ (.A1(net2157),
    .A2(net308),
    .B1(net348),
    .B2(_1442_),
    .X(_1474_));
 sky130_fd_sc_hd__a21oi_4 _3824_ (.A1(net1968),
    .A2(net356),
    .B1(net2158),
    .Y(_1475_));
 sky130_fd_sc_hd__nand2_1 _3825_ (.A(net379),
    .B(net2227),
    .Y(_1476_));
 sky130_fd_sc_hd__o21ai_4 _3826_ (.A1(net379),
    .A2(_1475_),
    .B1(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__inv_2 _3827_ (.A(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__and3_1 _3828_ (.A(net1968),
    .B(net367),
    .C(net350),
    .X(_1479_));
 sky130_fd_sc_hd__a221o_4 _3829_ (.A1(net2318),
    .A2(net305),
    .B1(net348),
    .B2(net307),
    .C1(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__nand2_1 _3830_ (.A(_1477_),
    .B(_1480_),
    .Y(_1481_));
 sky130_fd_sc_hd__or2_1 _3831_ (.A(_1477_),
    .B(_1480_),
    .X(_1482_));
 sky130_fd_sc_hd__and2b_1 _3832_ (.A_N(net437),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ),
    .X(_1483_));
 sky130_fd_sc_hd__a221o_1 _3833_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[30] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[30] ),
    .C1(_1483_),
    .X(_1484_));
 sky130_fd_sc_hd__mux2_1 _3834_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[30] ),
    .A1(_1484_),
    .S(net373),
    .X(_1485_));
 sky130_fd_sc_hd__and3_1 _3835_ (.A(net354),
    .B(net351),
    .C(net347),
    .X(_1486_));
 sky130_fd_sc_hd__a221o_2 _3836_ (.A1(net1992),
    .A2(net356),
    .B1(net308),
    .B2(net2281),
    .C1(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__mux2_2 _3837_ (.A0(net2259),
    .A1(_1487_),
    .S(net375),
    .X(_1488_));
 sky130_fd_sc_hd__and3_1 _3838_ (.A(net1992),
    .B(net367),
    .C(net350),
    .X(_1489_));
 sky130_fd_sc_hd__a221o_4 _3839_ (.A1(net2343),
    .A2(net305),
    .B1(_1485_),
    .B2(net307),
    .C1(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__nand2_1 _3840_ (.A(_1488_),
    .B(net2344),
    .Y(_1491_));
 sky130_fd_sc_hd__or2_1 _3841_ (.A(_1488_),
    .B(_1490_),
    .X(_1492_));
 sky130_fd_sc_hd__and2_1 _3842_ (.A(_1491_),
    .B(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__and2b_1 _3843_ (.A_N(net437),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[29] ),
    .X(_1494_));
 sky130_fd_sc_hd__a221o_1 _3844_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[29] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[29] ),
    .C1(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__mux2_1 _3845_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[29] ),
    .A1(_1495_),
    .S(net373),
    .X(_1496_));
 sky130_fd_sc_hd__a22o_1 _3846_ (.A1(net2236),
    .A2(net308),
    .B1(net346),
    .B2(_1442_),
    .X(_1497_));
 sky130_fd_sc_hd__a21oi_2 _3847_ (.A1(net2062),
    .A2(net356),
    .B1(net2237),
    .Y(_1498_));
 sky130_fd_sc_hd__nand2_1 _3848_ (.A(net379),
    .B(net2297),
    .Y(_1499_));
 sky130_fd_sc_hd__o21ai_4 _3849_ (.A1(net379),
    .A2(_1498_),
    .B1(net2298),
    .Y(_1500_));
 sky130_fd_sc_hd__inv_2 _3850_ (.A(_1500_),
    .Y(_1501_));
 sky130_fd_sc_hd__and3_1 _3851_ (.A(net2062),
    .B(net367),
    .C(net350),
    .X(_1502_));
 sky130_fd_sc_hd__a221o_4 _3852_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[29] ),
    .A2(net305),
    .B1(_1496_),
    .B2(net307),
    .C1(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__or2_1 _3853_ (.A(_1500_),
    .B(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__nand2_1 _3854_ (.A(_1500_),
    .B(_1503_),
    .Y(_1505_));
 sky130_fd_sc_hd__and2_1 _3855_ (.A(_1504_),
    .B(_1505_),
    .X(_1506_));
 sky130_fd_sc_hd__a2111o_2 _3856_ (.A1(_1481_),
    .A2(_1482_),
    .B1(_1493_),
    .C1(_1506_),
    .D1(_1469_),
    .X(_1507_));
 sky130_fd_sc_hd__and2b_1 _3857_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[17] ),
    .X(_1508_));
 sky130_fd_sc_hd__a221o_4 _3858_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[17] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[17] ),
    .C1(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__or2_2 _3859_ (.A(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[17] ),
    .B(net374),
    .X(_1510_));
 sky130_fd_sc_hd__o21ai_4 _3860_ (.A1(_1443_),
    .A2(_1509_),
    .B1(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__o21a_4 _3861_ (.A1(_1443_),
    .A2(_1509_),
    .B1(_1510_),
    .X(_1512_));
 sky130_fd_sc_hd__or3_1 _3862_ (.A(net355),
    .B(_1441_),
    .C(_1511_),
    .X(_1513_));
 sky130_fd_sc_hd__nand2_1 _3863_ (.A(net2067),
    .B(net355),
    .Y(_1514_));
 sky130_fd_sc_hd__or3b_1 _3864_ (.A(net355),
    .B(net351),
    .C_N(net2155),
    .X(_1515_));
 sky130_fd_sc_hd__a31o_1 _3865_ (.A1(_1513_),
    .A2(_1514_),
    .A3(_1515_),
    .B1(net380),
    .X(_1516_));
 sky130_fd_sc_hd__nand2_1 _3866_ (.A(net380),
    .B(net2209),
    .Y(_1517_));
 sky130_fd_sc_hd__nand2_2 _3867_ (.A(_1516_),
    .B(_1517_),
    .Y(_1518_));
 sky130_fd_sc_hd__and3_1 _3868_ (.A(net2067),
    .B(net366),
    .C(net349),
    .X(_1519_));
 sky130_fd_sc_hd__a221oi_4 _3869_ (.A1(net2323),
    .A2(net304),
    .B1(_1512_),
    .B2(net306),
    .C1(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__a221o_2 _3870_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ),
    .A2(net304),
    .B1(_1512_),
    .B2(net306),
    .C1(_1519_),
    .X(_1521_));
 sky130_fd_sc_hd__nand3_1 _3871_ (.A(_1516_),
    .B(_1517_),
    .C(_1520_),
    .Y(_1522_));
 sky130_fd_sc_hd__a21o_1 _3872_ (.A1(_1516_),
    .A2(_1517_),
    .B1(net2324),
    .X(_1523_));
 sky130_fd_sc_hd__and2b_1 _3873_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[19] ),
    .X(_1524_));
 sky130_fd_sc_hd__a221o_1 _3874_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[19] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[19] ),
    .C1(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__mux2_1 _3875_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[19] ),
    .A1(_1525_),
    .S(net374),
    .X(_1526_));
 sky130_fd_sc_hd__and3_1 _3876_ (.A(net353),
    .B(net351),
    .C(net345),
    .X(_1527_));
 sky130_fd_sc_hd__a221o_2 _3877_ (.A1(net767),
    .A2(net355),
    .B1(net309),
    .B2(net2220),
    .C1(_1527_),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_4 _3878_ (.A0(net2273),
    .A1(_1528_),
    .S(net375),
    .X(_1529_));
 sky130_fd_sc_hd__and3_1 _3879_ (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[19] ),
    .B(net366),
    .C(net349),
    .X(_1530_));
 sky130_fd_sc_hd__a221o_4 _3880_ (.A1(net2366),
    .A2(net304),
    .B1(net345),
    .B2(net306),
    .C1(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__or2_1 _3881_ (.A(_1529_),
    .B(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__nand2_1 _3882_ (.A(_1529_),
    .B(_1531_),
    .Y(_1533_));
 sky130_fd_sc_hd__and2_1 _3883_ (.A(_1532_),
    .B(_1533_),
    .X(_1534_));
 sky130_fd_sc_hd__and2b_1 _3884_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[16] ),
    .X(_1535_));
 sky130_fd_sc_hd__a221o_1 _3885_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[16] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[16] ),
    .C1(_1535_),
    .X(_1536_));
 sky130_fd_sc_hd__mux2_1 _3886_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[16] ),
    .A1(_1536_),
    .S(net373),
    .X(_1537_));
 sky130_fd_sc_hd__and3_1 _3887_ (.A(net354),
    .B(net351),
    .C(net344),
    .X(_1538_));
 sky130_fd_sc_hd__a221oi_4 _3888_ (.A1(net2122),
    .A2(net356),
    .B1(net308),
    .B2(net2313),
    .C1(_1538_),
    .Y(_1539_));
 sky130_fd_sc_hd__inv_2 _3889_ (.A(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__mux2_1 _3890_ (.A0(_1419_),
    .A1(_1539_),
    .S(net376),
    .X(_1541_));
 sky130_fd_sc_hd__mux2_1 _3891_ (.A0(net2252),
    .A1(_1540_),
    .S(net376),
    .X(_1542_));
 sky130_fd_sc_hd__and3_1 _3892_ (.A(net2122),
    .B(net367),
    .C(net350),
    .X(_1543_));
 sky130_fd_sc_hd__a221o_4 _3893_ (.A1(net2364),
    .A2(net305),
    .B1(_1537_),
    .B2(net307),
    .C1(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__nand2_1 _3894_ (.A(_1542_),
    .B(_1544_),
    .Y(_1545_));
 sky130_fd_sc_hd__or2_1 _3895_ (.A(_1542_),
    .B(_1544_),
    .X(_1546_));
 sky130_fd_sc_hd__and2_1 _3896_ (.A(_1545_),
    .B(_1546_),
    .X(_1547_));
 sky130_fd_sc_hd__and2b_1 _3897_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[18] ),
    .X(_1548_));
 sky130_fd_sc_hd__a221o_1 _3898_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[18] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[18] ),
    .C1(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__mux2_1 _3899_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[18] ),
    .A1(_1549_),
    .S(net373),
    .X(_1550_));
 sky130_fd_sc_hd__and3_1 _3900_ (.A(net353),
    .B(net351),
    .C(net343),
    .X(_1551_));
 sky130_fd_sc_hd__a221o_2 _3901_ (.A1(net1892),
    .A2(net355),
    .B1(net309),
    .B2(net2294),
    .C1(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__mux2_4 _3902_ (.A0(net2248),
    .A1(_1552_),
    .S(net375),
    .X(_1553_));
 sky130_fd_sc_hd__and3_1 _3903_ (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[18] ),
    .B(net366),
    .C(net349),
    .X(_1554_));
 sky130_fd_sc_hd__a221o_4 _3904_ (.A1(net2337),
    .A2(net304),
    .B1(net343),
    .B2(net306),
    .C1(_1554_),
    .X(_1555_));
 sky130_fd_sc_hd__nand2_1 _3905_ (.A(_1553_),
    .B(_1555_),
    .Y(_1556_));
 sky130_fd_sc_hd__or2_1 _3906_ (.A(_1553_),
    .B(_1555_),
    .X(_1557_));
 sky130_fd_sc_hd__xor2_1 _3907_ (.A(_1553_),
    .B(_1555_),
    .X(_1558_));
 sky130_fd_sc_hd__a2111o_2 _3908_ (.A1(_1522_),
    .A2(_1523_),
    .B1(_1534_),
    .C1(_1547_),
    .D1(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__and2b_1 _3909_ (.A_N(net437),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[21] ),
    .X(_1560_));
 sky130_fd_sc_hd__a221o_1 _3910_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[21] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[21] ),
    .C1(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__mux2_1 _3911_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[21] ),
    .A1(_1561_),
    .S(net373),
    .X(_1562_));
 sky130_fd_sc_hd__and3_1 _3912_ (.A(net354),
    .B(net351),
    .C(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__a221o_2 _3913_ (.A1(net1963),
    .A2(net356),
    .B1(net308),
    .B2(net2303),
    .C1(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__mux2_2 _3914_ (.A0(net2238),
    .A1(_1564_),
    .S(net375),
    .X(_1565_));
 sky130_fd_sc_hd__and3_1 _3915_ (.A(net1963),
    .B(net367),
    .C(net350),
    .X(_1566_));
 sky130_fd_sc_hd__a221o_4 _3916_ (.A1(net2341),
    .A2(net305),
    .B1(net342),
    .B2(net307),
    .C1(_1566_),
    .X(_1567_));
 sky130_fd_sc_hd__or2_1 _3917_ (.A(_1565_),
    .B(_1567_),
    .X(_1568_));
 sky130_fd_sc_hd__xor2_1 _3918_ (.A(_1565_),
    .B(_1567_),
    .X(_1569_));
 sky130_fd_sc_hd__and2b_1 _3919_ (.A_N(net437),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[22] ),
    .X(_1570_));
 sky130_fd_sc_hd__a221o_4 _3920_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[22] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[22] ),
    .C1(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__mux2_1 _3921_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[22] ),
    .A1(_1571_),
    .S(net374),
    .X(_1572_));
 sky130_fd_sc_hd__and3_1 _3922_ (.A(net353),
    .B(_1440_),
    .C(net341),
    .X(_1573_));
 sky130_fd_sc_hd__a221o_4 _3923_ (.A1(net1988),
    .A2(net357),
    .B1(net309),
    .B2(net2314),
    .C1(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__mux2_2 _3924_ (.A0(net2200),
    .A1(_1574_),
    .S(net375),
    .X(_1575_));
 sky130_fd_sc_hd__and3_1 _3925_ (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[22] ),
    .B(net366),
    .C(net349),
    .X(_1576_));
 sky130_fd_sc_hd__a221o_4 _3926_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ),
    .A2(net304),
    .B1(net341),
    .B2(net306),
    .C1(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__nand2_1 _3927_ (.A(_1575_),
    .B(_1577_),
    .Y(_1578_));
 sky130_fd_sc_hd__or2_1 _3928_ (.A(_1575_),
    .B(_1577_),
    .X(_1579_));
 sky130_fd_sc_hd__xor2_1 _3929_ (.A(_1575_),
    .B(_1577_),
    .X(_1580_));
 sky130_fd_sc_hd__or2_1 _3930_ (.A(_1569_),
    .B(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__and2b_1 _3931_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[20] ),
    .X(_1582_));
 sky130_fd_sc_hd__a221o_4 _3932_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[20] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[20] ),
    .C1(_1582_),
    .X(_1583_));
 sky130_fd_sc_hd__mux2_1 _3933_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[20] ),
    .A1(_1583_),
    .S(net373),
    .X(_1584_));
 sky130_fd_sc_hd__a22o_1 _3934_ (.A1(\U_DATAPATH.U_ID_EX.o_rs2_EX[20] ),
    .A2(net308),
    .B1(net340),
    .B2(_1442_),
    .X(_1585_));
 sky130_fd_sc_hd__a21oi_1 _3935_ (.A1(net2140),
    .A2(net356),
    .B1(_1585_),
    .Y(_1586_));
 sky130_fd_sc_hd__nand2_1 _3936_ (.A(net379),
    .B(net2160),
    .Y(_1587_));
 sky130_fd_sc_hd__o21ai_4 _3937_ (.A1(net379),
    .A2(net2141),
    .B1(_1587_),
    .Y(_1588_));
 sky130_fd_sc_hd__and3_1 _3938_ (.A(net2140),
    .B(net367),
    .C(net350),
    .X(_1589_));
 sky130_fd_sc_hd__a221o_4 _3939_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[20] ),
    .A2(net305),
    .B1(net340),
    .B2(net307),
    .C1(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__nand2_1 _3940_ (.A(_1588_),
    .B(_1590_),
    .Y(_1591_));
 sky130_fd_sc_hd__or2_1 _3941_ (.A(_1588_),
    .B(_1590_),
    .X(_1592_));
 sky130_fd_sc_hd__and2b_1 _3942_ (.A_N(net437),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[23] ),
    .X(_1593_));
 sky130_fd_sc_hd__a221o_1 _3943_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[23] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[23] ),
    .C1(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__mux2_1 _3944_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[23] ),
    .A1(_1594_),
    .S(net373),
    .X(_1595_));
 sky130_fd_sc_hd__a22o_1 _3945_ (.A1(net2267),
    .A2(net308),
    .B1(net339),
    .B2(_1442_),
    .X(_1596_));
 sky130_fd_sc_hd__a21oi_2 _3946_ (.A1(net2065),
    .A2(net356),
    .B1(net2268),
    .Y(_1597_));
 sky130_fd_sc_hd__nand2_1 _3947_ (.A(net379),
    .B(net2211),
    .Y(_1598_));
 sky130_fd_sc_hd__o21ai_4 _3948_ (.A1(net379),
    .A2(_1597_),
    .B1(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__and3_1 _3949_ (.A(net2065),
    .B(net367),
    .C(net350),
    .X(_1600_));
 sky130_fd_sc_hd__a221o_4 _3950_ (.A1(net2309),
    .A2(net305),
    .B1(_1595_),
    .B2(net307),
    .C1(_1600_),
    .X(_1601_));
 sky130_fd_sc_hd__or2_1 _3951_ (.A(_1599_),
    .B(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__xor2_1 _3952_ (.A(_1599_),
    .B(_1601_),
    .X(_1603_));
 sky130_fd_sc_hd__a211o_1 _3953_ (.A1(_1591_),
    .A2(_1592_),
    .B1(_1603_),
    .C1(_1581_),
    .X(_1604_));
 sky130_fd_sc_hd__and2b_1 _3954_ (.A_N(net437),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[25] ),
    .X(_1605_));
 sky130_fd_sc_hd__a221o_1 _3955_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[25] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[25] ),
    .C1(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__mux2_1 _3956_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[25] ),
    .A1(_1606_),
    .S(net373),
    .X(_1607_));
 sky130_fd_sc_hd__a22o_1 _3957_ (.A1(net2246),
    .A2(net308),
    .B1(net338),
    .B2(_1442_),
    .X(_1608_));
 sky130_fd_sc_hd__a21oi_4 _3958_ (.A1(net2153),
    .A2(net356),
    .B1(net2247),
    .Y(_1609_));
 sky130_fd_sc_hd__nand2_1 _3959_ (.A(net379),
    .B(net2216),
    .Y(_1610_));
 sky130_fd_sc_hd__o21ai_4 _3960_ (.A1(net379),
    .A2(_1609_),
    .B1(_1610_),
    .Y(_1611_));
 sky130_fd_sc_hd__inv_2 _3961_ (.A(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hd__and3_1 _3962_ (.A(net2153),
    .B(net367),
    .C(net350),
    .X(_1613_));
 sky130_fd_sc_hd__a221o_4 _3963_ (.A1(net2327),
    .A2(net305),
    .B1(net338),
    .B2(net307),
    .C1(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__or2_1 _3964_ (.A(_1611_),
    .B(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__xor2_1 _3965_ (.A(_1611_),
    .B(_1614_),
    .X(_1616_));
 sky130_fd_sc_hd__and2b_1 _3966_ (.A_N(net437),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[26] ),
    .X(_1617_));
 sky130_fd_sc_hd__a221o_1 _3967_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[26] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[26] ),
    .C1(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__mux2_1 _3968_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[26] ),
    .A1(_1618_),
    .S(net373),
    .X(_1619_));
 sky130_fd_sc_hd__and3_1 _3969_ (.A(net354),
    .B(net351),
    .C(net337),
    .X(_1620_));
 sky130_fd_sc_hd__a221o_2 _3970_ (.A1(net1993),
    .A2(net356),
    .B1(net308),
    .B2(net2276),
    .C1(_1620_),
    .X(_1621_));
 sky130_fd_sc_hd__mux2_2 _3971_ (.A0(net2305),
    .A1(_1621_),
    .S(net375),
    .X(_1622_));
 sky130_fd_sc_hd__and3_1 _3972_ (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[26] ),
    .B(net367),
    .C(net350),
    .X(_1623_));
 sky130_fd_sc_hd__a221o_4 _3973_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[26] ),
    .A2(net305),
    .B1(_1619_),
    .B2(net307),
    .C1(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__and2_1 _3974_ (.A(_1622_),
    .B(_1624_),
    .X(_1625_));
 sky130_fd_sc_hd__nor2_1 _3975_ (.A(_1622_),
    .B(_1624_),
    .Y(_1626_));
 sky130_fd_sc_hd__nor2_1 _3976_ (.A(_1625_),
    .B(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__and2b_1 _3977_ (.A_N(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[24] ),
    .X(_1628_));
 sky130_fd_sc_hd__a221o_1 _3978_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[24] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[24] ),
    .C1(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__mux2_2 _3979_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[24] ),
    .A1(_1629_),
    .S(net373),
    .X(_1630_));
 sky130_fd_sc_hd__a22o_1 _3980_ (.A1(net1156),
    .A2(net309),
    .B1(net336),
    .B2(_1442_),
    .X(_1631_));
 sky130_fd_sc_hd__a21oi_4 _3981_ (.A1(net863),
    .A2(net355),
    .B1(net1157),
    .Y(_1632_));
 sky130_fd_sc_hd__nand2_1 _3982_ (.A(net379),
    .B(net2123),
    .Y(_1633_));
 sky130_fd_sc_hd__o21ai_4 _3983_ (.A1(net379),
    .A2(_1632_),
    .B1(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__inv_2 _3984_ (.A(_1634_),
    .Y(_1635_));
 sky130_fd_sc_hd__and3_1 _3985_ (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[24] ),
    .B(net367),
    .C(net350),
    .X(_1636_));
 sky130_fd_sc_hd__a221o_4 _3986_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ),
    .A2(net305),
    .B1(net336),
    .B2(net307),
    .C1(_1636_),
    .X(_1637_));
 sky130_fd_sc_hd__and2_1 _3987_ (.A(_1634_),
    .B(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__nor2_1 _3988_ (.A(_1634_),
    .B(_1637_),
    .Y(_1639_));
 sky130_fd_sc_hd__nor2_1 _3989_ (.A(_1638_),
    .B(_1639_),
    .Y(_1640_));
 sky130_fd_sc_hd__and2b_1 _3990_ (.A_N(net437),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[27] ),
    .X(_1641_));
 sky130_fd_sc_hd__a221o_1 _3991_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[27] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[27] ),
    .C1(_1641_),
    .X(_1642_));
 sky130_fd_sc_hd__mux2_1 _3992_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[27] ),
    .A1(_1642_),
    .S(net373),
    .X(_1643_));
 sky130_fd_sc_hd__a22o_1 _3993_ (.A1(net2221),
    .A2(net308),
    .B1(net335),
    .B2(_1442_),
    .X(_1644_));
 sky130_fd_sc_hd__a21oi_2 _3994_ (.A1(net1991),
    .A2(net356),
    .B1(net2222),
    .Y(_1645_));
 sky130_fd_sc_hd__inv_2 _3995_ (.A(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__mux2_4 _3996_ (.A0(net2282),
    .A1(_1646_),
    .S(net375),
    .X(_1647_));
 sky130_fd_sc_hd__and3_1 _3997_ (.A(net1991),
    .B(net367),
    .C(net350),
    .X(_1648_));
 sky130_fd_sc_hd__a221o_4 _3998_ (.A1(net2328),
    .A2(net305),
    .B1(net335),
    .B2(net307),
    .C1(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__xor2_1 _3999_ (.A(_1647_),
    .B(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__or4_1 _4000_ (.A(_1616_),
    .B(_1627_),
    .C(_1640_),
    .D(_1650_),
    .X(_1651_));
 sky130_fd_sc_hd__or4_4 _4001_ (.A(_1507_),
    .B(_1559_),
    .C(_1604_),
    .D(_1651_),
    .X(_1652_));
 sky130_fd_sc_hd__and2b_1 _4002_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[3] ),
    .X(_1653_));
 sky130_fd_sc_hd__a221o_1 _4003_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[3] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[3] ),
    .C1(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__mux2_2 _4004_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[3] ),
    .A1(_1654_),
    .S(net374),
    .X(_1655_));
 sky130_fd_sc_hd__and3_1 _4005_ (.A(net353),
    .B(_1440_),
    .C(net334),
    .X(_1656_));
 sky130_fd_sc_hd__a221oi_4 _4006_ (.A1(\U_DATAPATH.U_EX_MEM.o_alu_result_M[3] ),
    .A2(net355),
    .B1(net309),
    .B2(net2120),
    .C1(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__nand2_2 _4007_ (.A(net380),
    .B(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ),
    .Y(_1658_));
 sky130_fd_sc_hd__o21a_4 _4008_ (.A1(net380),
    .A2(_1657_),
    .B1(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__o21ai_4 _4009_ (.A1(net380),
    .A2(_1657_),
    .B1(_1658_),
    .Y(_1660_));
 sky130_fd_sc_hd__and3_1 _4010_ (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[3] ),
    .B(net366),
    .C(net349),
    .X(_1661_));
 sky130_fd_sc_hd__a221o_4 _4011_ (.A1(net2365),
    .A2(net304),
    .B1(net334),
    .B2(net306),
    .C1(_1661_),
    .X(_1662_));
 sky130_fd_sc_hd__or2_1 _4012_ (.A(net211),
    .B(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__xnor2_1 _4013_ (.A(net211),
    .B(_1662_),
    .Y(_1664_));
 sky130_fd_sc_hd__and2b_1 _4014_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[2] ),
    .X(_1665_));
 sky130_fd_sc_hd__a221o_1 _4015_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[2] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[2] ),
    .C1(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__mux2_2 _4016_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[2] ),
    .A1(_1666_),
    .S(net374),
    .X(_1667_));
 sky130_fd_sc_hd__and3_1 _4017_ (.A(net353),
    .B(_1440_),
    .C(net333),
    .X(_1668_));
 sky130_fd_sc_hd__a221o_4 _4018_ (.A1(net1780),
    .A2(net357),
    .B1(net309),
    .B2(net2317),
    .C1(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__and2_1 _4019_ (.A(net380),
    .B(net2333),
    .X(_1670_));
 sky130_fd_sc_hd__a21oi_1 _4020_ (.A1(net376),
    .A2(_1669_),
    .B1(_1670_),
    .Y(_1671_));
 sky130_fd_sc_hd__a21o_1 _4021_ (.A1(net376),
    .A2(_1669_),
    .B1(_1670_),
    .X(_1672_));
 sky130_fd_sc_hd__and3_1 _4022_ (.A(net1780),
    .B(net366),
    .C(net349),
    .X(_1673_));
 sky130_fd_sc_hd__a221o_4 _4023_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[2] ),
    .A2(net304),
    .B1(net333),
    .B2(net306),
    .C1(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__nand2_1 _4024_ (.A(_1672_),
    .B(_1674_),
    .Y(_1675_));
 sky130_fd_sc_hd__xnor2_1 _4025_ (.A(net204),
    .B(_1674_),
    .Y(_1676_));
 sky130_fd_sc_hd__nand2_1 _4026_ (.A(_1664_),
    .B(_1676_),
    .Y(_1677_));
 sky130_fd_sc_hd__a22o_1 _4027_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[1] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[1] ),
    .X(_1678_));
 sky130_fd_sc_hd__a21o_2 _4028_ (.A1(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[1] ),
    .A2(_1443_),
    .B1(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__and3_1 _4029_ (.A(net353),
    .B(net351),
    .C(net332),
    .X(_1680_));
 sky130_fd_sc_hd__nor2_1 _4030_ (.A(_1420_),
    .B(net353),
    .Y(_1681_));
 sky130_fd_sc_hd__and3_2 _4031_ (.A(net2330),
    .B(net353),
    .C(_1441_),
    .X(_1682_));
 sky130_fd_sc_hd__o31a_1 _4032_ (.A1(_1680_),
    .A2(_1681_),
    .A3(_1682_),
    .B1(net376),
    .X(_1683_));
 sky130_fd_sc_hd__nand2_1 _4033_ (.A(net380),
    .B(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[1] ),
    .Y(_1684_));
 sky130_fd_sc_hd__inv_2 _4034_ (.A(_1684_),
    .Y(_1685_));
 sky130_fd_sc_hd__nor2_2 _4035_ (.A(_1683_),
    .B(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hd__or2_1 _4036_ (.A(_1683_),
    .B(_1685_),
    .X(_1687_));
 sky130_fd_sc_hd__and3_1 _4037_ (.A(net1507),
    .B(net366),
    .C(net349),
    .X(_1688_));
 sky130_fd_sc_hd__a221o_4 _4038_ (.A1(net2363),
    .A2(net304),
    .B1(net332),
    .B2(net306),
    .C1(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__inv_2 _4039_ (.A(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__or2_1 _4040_ (.A(net199),
    .B(_1689_),
    .X(_1691_));
 sky130_fd_sc_hd__nand2_1 _4041_ (.A(net199),
    .B(_1689_),
    .Y(_1692_));
 sky130_fd_sc_hd__and2_1 _4042_ (.A(_1691_),
    .B(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__a22o_1 _4043_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[0] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[0] ),
    .X(_1694_));
 sky130_fd_sc_hd__a21o_1 _4044_ (.A1(net2045),
    .A2(_1443_),
    .B1(_1694_),
    .X(_1695_));
 sky130_fd_sc_hd__and3_1 _4045_ (.A(net353),
    .B(net351),
    .C(net331),
    .X(_1696_));
 sky130_fd_sc_hd__a221o_1 _4046_ (.A1(net2133),
    .A2(net355),
    .B1(net309),
    .B2(net2326),
    .C1(_1696_),
    .X(_1697_));
 sky130_fd_sc_hd__mux2_2 _4047_ (.A0(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[0] ),
    .A1(_1697_),
    .S(net376),
    .X(_1698_));
 sky130_fd_sc_hd__inv_2 _4048_ (.A(net192),
    .Y(_1699_));
 sky130_fd_sc_hd__and3_1 _4049_ (.A(net2133),
    .B(net366),
    .C(net349),
    .X(_1700_));
 sky130_fd_sc_hd__a221o_4 _4050_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ),
    .A2(net304),
    .B1(net331),
    .B2(net306),
    .C1(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__inv_2 _4051_ (.A(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hd__nand2_1 _4052_ (.A(net195),
    .B(_1701_),
    .Y(_1703_));
 sky130_fd_sc_hd__or2_1 _4053_ (.A(net195),
    .B(_1701_),
    .X(_1704_));
 sky130_fd_sc_hd__and2b_1 _4054_ (.A_N(net437),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[7] ),
    .X(_1705_));
 sky130_fd_sc_hd__a221o_4 _4055_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[7] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[7] ),
    .C1(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__mux2_1 _4056_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[7] ),
    .A1(_1706_),
    .S(net373),
    .X(_1707_));
 sky130_fd_sc_hd__and3_1 _4057_ (.A(net354),
    .B(net351),
    .C(net330),
    .X(_1708_));
 sky130_fd_sc_hd__a221o_4 _4058_ (.A1(net2054),
    .A2(net356),
    .B1(net308),
    .B2(net2196),
    .C1(_1708_),
    .X(_1709_));
 sky130_fd_sc_hd__mux2_4 _4059_ (.A0(net2184),
    .A1(_1709_),
    .S(net375),
    .X(_1710_));
 sky130_fd_sc_hd__and3_1 _4060_ (.A(net2054),
    .B(net367),
    .C(net350),
    .X(_1711_));
 sky130_fd_sc_hd__a221o_4 _4061_ (.A1(net2357),
    .A2(net305),
    .B1(_1707_),
    .B2(net307),
    .C1(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__xor2_1 _4062_ (.A(_1710_),
    .B(_1712_),
    .X(_1713_));
 sky130_fd_sc_hd__and2b_1 _4063_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[4] ),
    .X(_1714_));
 sky130_fd_sc_hd__a221o_2 _4064_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[4] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[4] ),
    .C1(_1714_),
    .X(_1715_));
 sky130_fd_sc_hd__mux2_1 _4065_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[4] ),
    .A1(_1715_),
    .S(net374),
    .X(_1716_));
 sky130_fd_sc_hd__and3_1 _4066_ (.A(net354),
    .B(net352),
    .C(net329),
    .X(_1717_));
 sky130_fd_sc_hd__a221o_4 _4067_ (.A1(net2127),
    .A2(net355),
    .B1(net309),
    .B2(net2231),
    .C1(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__and2_1 _4068_ (.A(net380),
    .B(net2295),
    .X(_1719_));
 sky130_fd_sc_hd__a21oi_1 _4069_ (.A1(net375),
    .A2(_1718_),
    .B1(_1719_),
    .Y(_1720_));
 sky130_fd_sc_hd__a21o_2 _4070_ (.A1(net375),
    .A2(_1718_),
    .B1(_1719_),
    .X(_1721_));
 sky130_fd_sc_hd__and3_1 _4071_ (.A(net2127),
    .B(_1453_),
    .C(_1457_),
    .X(_1722_));
 sky130_fd_sc_hd__a221o_4 _4072_ (.A1(net2371),
    .A2(net304),
    .B1(net329),
    .B2(net306),
    .C1(_1722_),
    .X(_1723_));
 sky130_fd_sc_hd__nand2_1 _4073_ (.A(net188),
    .B(_1723_),
    .Y(_1724_));
 sky130_fd_sc_hd__or2_1 _4074_ (.A(net188),
    .B(_1723_),
    .X(_1725_));
 sky130_fd_sc_hd__and2b_1 _4075_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[6] ),
    .X(_1726_));
 sky130_fd_sc_hd__a221o_1 _4076_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[6] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[6] ),
    .C1(_1726_),
    .X(_1727_));
 sky130_fd_sc_hd__mux2_1 _4077_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[6] ),
    .A1(_1727_),
    .S(net374),
    .X(_1728_));
 sky130_fd_sc_hd__and3_1 _4078_ (.A(net353),
    .B(net352),
    .C(net328),
    .X(_1729_));
 sky130_fd_sc_hd__a221o_1 _4079_ (.A1(net2159),
    .A2(net355),
    .B1(net309),
    .B2(net2175),
    .C1(_1729_),
    .X(_1730_));
 sky130_fd_sc_hd__mux2_2 _4080_ (.A0(net2177),
    .A1(_1730_),
    .S(net376),
    .X(_1731_));
 sky130_fd_sc_hd__and3_1 _4081_ (.A(net2159),
    .B(net366),
    .C(net349),
    .X(_1732_));
 sky130_fd_sc_hd__a221o_4 _4082_ (.A1(net2331),
    .A2(net304),
    .B1(net328),
    .B2(net306),
    .C1(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__nand2_1 _4083_ (.A(_1731_),
    .B(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__or2_1 _4084_ (.A(_1731_),
    .B(_1733_),
    .X(_1735_));
 sky130_fd_sc_hd__xor2_1 _4085_ (.A(_1731_),
    .B(_1733_),
    .X(_1736_));
 sky130_fd_sc_hd__and2b_1 _4086_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[5] ),
    .X(_1737_));
 sky130_fd_sc_hd__a221o_2 _4087_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[5] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[5] ),
    .C1(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__or2_2 _4088_ (.A(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[5] ),
    .B(net374),
    .X(_1739_));
 sky130_fd_sc_hd__o21ai_4 _4089_ (.A1(_1443_),
    .A2(_1738_),
    .B1(_1739_),
    .Y(_1740_));
 sky130_fd_sc_hd__o21a_4 _4090_ (.A1(_1443_),
    .A2(_1738_),
    .B1(_1739_),
    .X(_1741_));
 sky130_fd_sc_hd__and3_1 _4091_ (.A(net353),
    .B(net352),
    .C(_1741_),
    .X(_1742_));
 sky130_fd_sc_hd__and2_1 _4092_ (.A(net2035),
    .B(net355),
    .X(_1743_));
 sky130_fd_sc_hd__and3_1 _4093_ (.A(net2272),
    .B(net353),
    .C(_1441_),
    .X(_1744_));
 sky130_fd_sc_hd__o31a_2 _4094_ (.A1(_1742_),
    .A2(_1743_),
    .A3(_1744_),
    .B1(net375),
    .X(_1745_));
 sky130_fd_sc_hd__and2_1 _4095_ (.A(net380),
    .B(net2191),
    .X(_1746_));
 sky130_fd_sc_hd__or2_1 _4096_ (.A(_1745_),
    .B(_1746_),
    .X(_1747_));
 sky130_fd_sc_hd__and3_1 _4097_ (.A(net2035),
    .B(net366),
    .C(net349),
    .X(_1748_));
 sky130_fd_sc_hd__a221o_4 _4098_ (.A1(net2321),
    .A2(net304),
    .B1(_1741_),
    .B2(net306),
    .C1(_1748_),
    .X(_1749_));
 sky130_fd_sc_hd__or3_1 _4099_ (.A(_1745_),
    .B(_1746_),
    .C(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__o21ai_1 _4100_ (.A1(_1745_),
    .A2(_1746_),
    .B1(_1749_),
    .Y(_1751_));
 sky130_fd_sc_hd__and2_1 _4101_ (.A(_1750_),
    .B(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__a2111o_1 _4102_ (.A1(_1724_),
    .A2(_1725_),
    .B1(_1736_),
    .C1(_1752_),
    .D1(_1713_),
    .X(_1753_));
 sky130_fd_sc_hd__a2111o_1 _4103_ (.A1(_1703_),
    .A2(_1704_),
    .B1(_1753_),
    .C1(_1693_),
    .D1(_1677_),
    .X(_1754_));
 sky130_fd_sc_hd__and2b_1 _4104_ (.A_N(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[9] ),
    .X(_1755_));
 sky130_fd_sc_hd__a221o_1 _4105_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[9] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[9] ),
    .C1(_1755_),
    .X(_1756_));
 sky130_fd_sc_hd__mux2_1 _4106_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[9] ),
    .A1(_1756_),
    .S(net374),
    .X(_1757_));
 sky130_fd_sc_hd__and3_1 _4107_ (.A(net353),
    .B(net352),
    .C(net327),
    .X(_1758_));
 sky130_fd_sc_hd__a221o_4 _4108_ (.A1(net1919),
    .A2(net355),
    .B1(net309),
    .B2(net2245),
    .C1(_1758_),
    .X(_1759_));
 sky130_fd_sc_hd__mux2_2 _4109_ (.A0(net2274),
    .A1(_1759_),
    .S(net375),
    .X(_1760_));
 sky130_fd_sc_hd__and3_1 _4110_ (.A(net1919),
    .B(net366),
    .C(net349),
    .X(_1761_));
 sky130_fd_sc_hd__a221o_4 _4111_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ),
    .A2(net304),
    .B1(net327),
    .B2(net306),
    .C1(_1761_),
    .X(_1762_));
 sky130_fd_sc_hd__or2_1 _4112_ (.A(_1760_),
    .B(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__xor2_1 _4113_ (.A(_1760_),
    .B(_1762_),
    .X(_1764_));
 sky130_fd_sc_hd__and2b_1 _4114_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[10] ),
    .X(_1765_));
 sky130_fd_sc_hd__a221o_1 _4115_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[10] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[10] ),
    .C1(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__mux2_1 _4116_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[10] ),
    .A1(_1766_),
    .S(net373),
    .X(_1767_));
 sky130_fd_sc_hd__and3_1 _4117_ (.A(net354),
    .B(net351),
    .C(net326),
    .X(_1768_));
 sky130_fd_sc_hd__a221o_4 _4118_ (.A1(net2066),
    .A2(net356),
    .B1(net308),
    .B2(net2173),
    .C1(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__mux2_2 _4119_ (.A0(net2270),
    .A1(_1769_),
    .S(net375),
    .X(_1770_));
 sky130_fd_sc_hd__and3_1 _4120_ (.A(net2066),
    .B(net367),
    .C(net350),
    .X(_1771_));
 sky130_fd_sc_hd__a221o_4 _4121_ (.A1(net2339),
    .A2(net305),
    .B1(net326),
    .B2(net307),
    .C1(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__nand2_1 _4122_ (.A(_1770_),
    .B(_1772_),
    .Y(_1773_));
 sky130_fd_sc_hd__xor2_1 _4123_ (.A(_1770_),
    .B(_1772_),
    .X(_1774_));
 sky130_fd_sc_hd__and2b_1 _4124_ (.A_N(net437),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[8] ),
    .X(_1775_));
 sky130_fd_sc_hd__a221o_1 _4125_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[8] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[8] ),
    .C1(_1775_),
    .X(_1776_));
 sky130_fd_sc_hd__mux2_1 _4126_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[8] ),
    .A1(_1776_),
    .S(net373),
    .X(_1777_));
 sky130_fd_sc_hd__a22o_1 _4127_ (.A1(net2164),
    .A2(net308),
    .B1(net325),
    .B2(_1442_),
    .X(_1778_));
 sky130_fd_sc_hd__a21oi_4 _4128_ (.A1(net2139),
    .A2(net356),
    .B1(net2165),
    .Y(_1779_));
 sky130_fd_sc_hd__nand2_1 _4129_ (.A(net379),
    .B(net2301),
    .Y(_1780_));
 sky130_fd_sc_hd__o21ai_4 _4130_ (.A1(net379),
    .A2(_1779_),
    .B1(_1780_),
    .Y(_1781_));
 sky130_fd_sc_hd__and3_1 _4131_ (.A(net2139),
    .B(net367),
    .C(net350),
    .X(_1782_));
 sky130_fd_sc_hd__a221o_4 _4132_ (.A1(net2319),
    .A2(net305),
    .B1(_1777_),
    .B2(net307),
    .C1(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__nand2_1 _4133_ (.A(_1781_),
    .B(net2320),
    .Y(_1784_));
 sky130_fd_sc_hd__or2_1 _4134_ (.A(_1781_),
    .B(_1783_),
    .X(_1785_));
 sky130_fd_sc_hd__and2b_1 _4135_ (.A_N(net437),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[11] ),
    .X(_1786_));
 sky130_fd_sc_hd__a221o_1 _4136_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[11] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[11] ),
    .C1(_1786_),
    .X(_1787_));
 sky130_fd_sc_hd__mux2_1 _4137_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[11] ),
    .A1(_1787_),
    .S(net373),
    .X(_1788_));
 sky130_fd_sc_hd__and3_1 _4138_ (.A(net354),
    .B(net351),
    .C(net324),
    .X(_1789_));
 sky130_fd_sc_hd__a221o_2 _4139_ (.A1(net2009),
    .A2(net356),
    .B1(net308),
    .B2(net2205),
    .C1(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__mux2_4 _4140_ (.A0(net2359),
    .A1(_1790_),
    .S(net375),
    .X(_1791_));
 sky130_fd_sc_hd__and3_1 _4141_ (.A(net2009),
    .B(net367),
    .C(net350),
    .X(_1792_));
 sky130_fd_sc_hd__a221o_4 _4142_ (.A1(net2361),
    .A2(net305),
    .B1(_1788_),
    .B2(net307),
    .C1(_1792_),
    .X(_1793_));
 sky130_fd_sc_hd__or2_1 _4143_ (.A(_1791_),
    .B(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__xor2_1 _4144_ (.A(_1791_),
    .B(_1793_),
    .X(_1795_));
 sky130_fd_sc_hd__or3_1 _4145_ (.A(_1764_),
    .B(_1774_),
    .C(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__a21o_1 _4146_ (.A1(_1784_),
    .A2(_1785_),
    .B1(_1796_),
    .X(_1797_));
 sky130_fd_sc_hd__and2b_1 _4147_ (.A_N(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[13] ),
    .X(_1798_));
 sky130_fd_sc_hd__a221o_1 _4148_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[13] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[13] ),
    .C1(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__mux2_1 _4149_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[13] ),
    .A1(_1799_),
    .S(net374),
    .X(_1800_));
 sky130_fd_sc_hd__and3_1 _4150_ (.A(net353),
    .B(net351),
    .C(net323),
    .X(_1801_));
 sky130_fd_sc_hd__a221o_4 _4151_ (.A1(net2091),
    .A2(net357),
    .B1(net309),
    .B2(net2285),
    .C1(_1801_),
    .X(_1802_));
 sky130_fd_sc_hd__mux2_2 _4152_ (.A0(net2286),
    .A1(_1802_),
    .S(net376),
    .X(_1803_));
 sky130_fd_sc_hd__inv_2 _4153_ (.A(_1803_),
    .Y(_1804_));
 sky130_fd_sc_hd__and3_1 _4154_ (.A(net2091),
    .B(net366),
    .C(net349),
    .X(_1805_));
 sky130_fd_sc_hd__a221o_4 _4155_ (.A1(net2336),
    .A2(net304),
    .B1(net323),
    .B2(net306),
    .C1(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__xor2_1 _4156_ (.A(_1803_),
    .B(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__and2b_1 _4157_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[14] ),
    .X(_1808_));
 sky130_fd_sc_hd__a221o_1 _4158_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[14] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[14] ),
    .C1(_1808_),
    .X(_1809_));
 sky130_fd_sc_hd__mux2_2 _4159_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[14] ),
    .A1(_1809_),
    .S(net374),
    .X(_1810_));
 sky130_fd_sc_hd__and3_1 _4160_ (.A(net353),
    .B(net351),
    .C(net322),
    .X(_1811_));
 sky130_fd_sc_hd__a221o_2 _4161_ (.A1(net2025),
    .A2(net355),
    .B1(net308),
    .B2(net2292),
    .C1(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__mux2_2 _4162_ (.A0(net2241),
    .A1(_1812_),
    .S(net375),
    .X(_1813_));
 sky130_fd_sc_hd__and3_1 _4163_ (.A(net2025),
    .B(net366),
    .C(net349),
    .X(_1814_));
 sky130_fd_sc_hd__a221o_4 _4164_ (.A1(net2353),
    .A2(_1466_),
    .B1(net322),
    .B2(net306),
    .C1(_1814_),
    .X(_1815_));
 sky130_fd_sc_hd__and2_1 _4165_ (.A(_1813_),
    .B(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__nor2_1 _4166_ (.A(_1813_),
    .B(_1815_),
    .Y(_1817_));
 sky130_fd_sc_hd__nor2_1 _4167_ (.A(_1816_),
    .B(_1817_),
    .Y(_1818_));
 sky130_fd_sc_hd__and2b_1 _4168_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[12] ),
    .X(_1819_));
 sky130_fd_sc_hd__a221o_2 _4169_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[12] ),
    .A2(net371),
    .B1(net368),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[12] ),
    .C1(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__mux2_1 _4170_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[12] ),
    .A1(_1820_),
    .S(net374),
    .X(_1821_));
 sky130_fd_sc_hd__a22o_1 _4171_ (.A1(net2084),
    .A2(net309),
    .B1(net321),
    .B2(_1442_),
    .X(_1822_));
 sky130_fd_sc_hd__a21oi_4 _4172_ (.A1(net1822),
    .A2(net355),
    .B1(net2085),
    .Y(_1823_));
 sky130_fd_sc_hd__nand2_1 _4173_ (.A(net380),
    .B(net2223),
    .Y(_1824_));
 sky130_fd_sc_hd__o21ai_4 _4174_ (.A1(net380),
    .A2(_1823_),
    .B1(_1824_),
    .Y(_1825_));
 sky130_fd_sc_hd__inv_2 _4175_ (.A(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__and3_1 _4176_ (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[12] ),
    .B(net366),
    .C(net349),
    .X(_1827_));
 sky130_fd_sc_hd__a221o_4 _4177_ (.A1(net2349),
    .A2(net304),
    .B1(net321),
    .B2(net306),
    .C1(_1827_),
    .X(_1828_));
 sky130_fd_sc_hd__and2_1 _4178_ (.A(_1825_),
    .B(net2350),
    .X(_1829_));
 sky130_fd_sc_hd__nor2_1 _4179_ (.A(_1825_),
    .B(_1828_),
    .Y(_1830_));
 sky130_fd_sc_hd__nor2_1 _4180_ (.A(_1829_),
    .B(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__and2b_1 _4181_ (.A_N(net438),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[15] ),
    .X(_1832_));
 sky130_fd_sc_hd__a221o_1 _4182_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[15] ),
    .A2(net372),
    .B1(net369),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[15] ),
    .C1(_1832_),
    .X(_1833_));
 sky130_fd_sc_hd__mux2_1 _4183_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[15] ),
    .A1(_1833_),
    .S(net374),
    .X(_1834_));
 sky130_fd_sc_hd__and3_1 _4184_ (.A(net353),
    .B(net351),
    .C(net320),
    .X(_1835_));
 sky130_fd_sc_hd__a221o_1 _4185_ (.A1(net1709),
    .A2(net355),
    .B1(net309),
    .B2(net2142),
    .C1(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__mux2_2 _4186_ (.A0(net2279),
    .A1(_1836_),
    .S(net375),
    .X(_1837_));
 sky130_fd_sc_hd__and3_1 _4187_ (.A(net1709),
    .B(_1453_),
    .C(_1457_),
    .X(_1838_));
 sky130_fd_sc_hd__a221o_4 _4188_ (.A1(net2345),
    .A2(net304),
    .B1(_1834_),
    .B2(_1464_),
    .C1(_1838_),
    .X(_1839_));
 sky130_fd_sc_hd__or2_1 _4189_ (.A(_1837_),
    .B(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__nand2_1 _4190_ (.A(_1837_),
    .B(_1839_),
    .Y(_1841_));
 sky130_fd_sc_hd__and2_1 _4191_ (.A(_1840_),
    .B(_1841_),
    .X(_1842_));
 sky130_fd_sc_hd__or4_2 _4192_ (.A(_1807_),
    .B(_1818_),
    .C(_1831_),
    .D(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__or4_4 _4193_ (.A(_1652_),
    .B(_1754_),
    .C(_1797_),
    .D(_1843_),
    .X(_1844_));
 sky130_fd_sc_hd__nand2b_1 _4194_ (.A_N(_1733_),
    .B(_1731_),
    .Y(_1845_));
 sky130_fd_sc_hd__nand2b_1 _4195_ (.A_N(_1749_),
    .B(_1747_),
    .Y(_1846_));
 sky130_fd_sc_hd__a211o_1 _4196_ (.A1(_1750_),
    .A2(_1751_),
    .B1(net191),
    .C1(_1723_),
    .X(_1847_));
 sky130_fd_sc_hd__a21o_1 _4197_ (.A1(_1846_),
    .A2(_1847_),
    .B1(_1736_),
    .X(_1848_));
 sky130_fd_sc_hd__a21o_1 _4198_ (.A1(_1845_),
    .A2(_1848_),
    .B1(_1713_),
    .X(_1849_));
 sky130_fd_sc_hd__nand2b_1 _4199_ (.A_N(_1712_),
    .B(_1710_),
    .Y(_1850_));
 sky130_fd_sc_hd__o21a_1 _4200_ (.A1(net196),
    .A2(_1702_),
    .B1(net199),
    .X(_1851_));
 sky130_fd_sc_hd__or3_2 _4201_ (.A(net199),
    .B(net196),
    .C(_1702_),
    .X(_1852_));
 sky130_fd_sc_hd__o2111ai_1 _4202_ (.A1(_1690_),
    .A2(_1851_),
    .B1(_1852_),
    .C1(_1676_),
    .D1(_1664_),
    .Y(_1853_));
 sky130_fd_sc_hd__or2_1 _4203_ (.A(_1659_),
    .B(_1662_),
    .X(_1854_));
 sky130_fd_sc_hd__or3b_1 _4204_ (.A(_1674_),
    .B(net207),
    .C_N(_1664_),
    .X(_1855_));
 sky130_fd_sc_hd__a31o_1 _4205_ (.A1(_1853_),
    .A2(_1854_),
    .A3(_1855_),
    .B1(_1753_),
    .X(_1856_));
 sky130_fd_sc_hd__a31o_1 _4206_ (.A1(_1849_),
    .A2(_1850_),
    .A3(_1856_),
    .B1(_1797_),
    .X(_1857_));
 sky130_fd_sc_hd__nand2b_1 _4207_ (.A_N(_1772_),
    .B(_1770_),
    .Y(_1858_));
 sky130_fd_sc_hd__nand2b_1 _4208_ (.A_N(_1762_),
    .B(_1760_),
    .Y(_1859_));
 sky130_fd_sc_hd__or3b_1 _4209_ (.A(_1764_),
    .B(_1783_),
    .C_N(_1781_),
    .X(_1860_));
 sky130_fd_sc_hd__a21o_1 _4210_ (.A1(_1859_),
    .A2(_1860_),
    .B1(_1774_),
    .X(_1861_));
 sky130_fd_sc_hd__a21o_1 _4211_ (.A1(_1858_),
    .A2(_1861_),
    .B1(_1795_),
    .X(_1862_));
 sky130_fd_sc_hd__nand2b_1 _4212_ (.A_N(_1793_),
    .B(_1791_),
    .Y(_1863_));
 sky130_fd_sc_hd__a31o_1 _4213_ (.A1(_1857_),
    .A2(_1862_),
    .A3(_1863_),
    .B1(_1843_),
    .X(_1864_));
 sky130_fd_sc_hd__nand2b_1 _4214_ (.A_N(_1815_),
    .B(_1813_),
    .Y(_1865_));
 sky130_fd_sc_hd__o32a_1 _4215_ (.A1(_1807_),
    .A2(_1826_),
    .A3(_1828_),
    .B1(_1806_),
    .B2(_1804_),
    .X(_1866_));
 sky130_fd_sc_hd__o21a_1 _4216_ (.A1(_1818_),
    .A2(_1866_),
    .B1(_1865_),
    .X(_1867_));
 sky130_fd_sc_hd__or2_1 _4217_ (.A(_1842_),
    .B(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__nand2b_1 _4218_ (.A_N(_1839_),
    .B(_1837_),
    .Y(_1869_));
 sky130_fd_sc_hd__a31oi_1 _4219_ (.A1(_1864_),
    .A2(_1868_),
    .A3(_1869_),
    .B1(_1652_),
    .Y(_1870_));
 sky130_fd_sc_hd__nand2_1 _4220_ (.A(_1451_),
    .B(_1468_),
    .Y(_1871_));
 sky130_fd_sc_hd__nand2b_1 _4221_ (.A_N(_1490_),
    .B(_1488_),
    .Y(_1872_));
 sky130_fd_sc_hd__o32a_1 _4222_ (.A1(_1478_),
    .A2(_1480_),
    .A3(_1506_),
    .B1(_1503_),
    .B2(_1501_),
    .X(_1873_));
 sky130_fd_sc_hd__o21a_1 _4223_ (.A1(_1493_),
    .A2(_1873_),
    .B1(_1872_),
    .X(_1874_));
 sky130_fd_sc_hd__o21ai_2 _4224_ (.A1(_1469_),
    .A2(_1874_),
    .B1(_1871_),
    .Y(_1875_));
 sky130_fd_sc_hd__nand2b_1 _4225_ (.A_N(_1531_),
    .B(_1529_),
    .Y(_1876_));
 sky130_fd_sc_hd__nand2b_1 _4226_ (.A_N(_1555_),
    .B(_1553_),
    .Y(_1877_));
 sky130_fd_sc_hd__and2_1 _4227_ (.A(_1518_),
    .B(_1520_),
    .X(_1878_));
 sky130_fd_sc_hd__a211oi_1 _4228_ (.A1(_1522_),
    .A2(_1523_),
    .B1(_1541_),
    .C1(_1544_),
    .Y(_1879_));
 sky130_fd_sc_hd__o21bai_1 _4229_ (.A1(_1878_),
    .A2(_1879_),
    .B1_N(_1558_),
    .Y(_1880_));
 sky130_fd_sc_hd__a21o_1 _4230_ (.A1(_1877_),
    .A2(_1880_),
    .B1(_1534_),
    .X(_1881_));
 sky130_fd_sc_hd__a21o_1 _4231_ (.A1(_1876_),
    .A2(_1881_),
    .B1(_1604_),
    .X(_1882_));
 sky130_fd_sc_hd__nand2b_1 _4232_ (.A_N(_1577_),
    .B(_1575_),
    .Y(_1883_));
 sky130_fd_sc_hd__nand2b_1 _4233_ (.A_N(_1567_),
    .B(_1565_),
    .Y(_1884_));
 sky130_fd_sc_hd__or3b_1 _4234_ (.A(_1569_),
    .B(_1590_),
    .C_N(_1588_),
    .X(_1885_));
 sky130_fd_sc_hd__a21o_1 _4235_ (.A1(_1884_),
    .A2(_1885_),
    .B1(_1580_),
    .X(_1886_));
 sky130_fd_sc_hd__a21o_1 _4236_ (.A1(_1883_),
    .A2(_1886_),
    .B1(_1603_),
    .X(_1887_));
 sky130_fd_sc_hd__nand2b_1 _4237_ (.A_N(_1601_),
    .B(_1599_),
    .Y(_1888_));
 sky130_fd_sc_hd__a31o_1 _4238_ (.A1(_1882_),
    .A2(_1887_),
    .A3(_1888_),
    .B1(_1651_),
    .X(_1889_));
 sky130_fd_sc_hd__nand2b_1 _4239_ (.A_N(_1624_),
    .B(_1622_),
    .Y(_1890_));
 sky130_fd_sc_hd__o32a_1 _4240_ (.A1(_1616_),
    .A2(_1635_),
    .A3(_1637_),
    .B1(_1614_),
    .B2(_1612_),
    .X(_1891_));
 sky130_fd_sc_hd__o21a_1 _4241_ (.A1(_1627_),
    .A2(_1891_),
    .B1(_1890_),
    .X(_1892_));
 sky130_fd_sc_hd__or2_1 _4242_ (.A(_1650_),
    .B(_1892_),
    .X(_1893_));
 sky130_fd_sc_hd__nand2b_1 _4243_ (.A_N(_1649_),
    .B(_1647_),
    .Y(_1894_));
 sky130_fd_sc_hd__a31oi_4 _4244_ (.A1(_1889_),
    .A2(_1893_),
    .A3(_1894_),
    .B1(_1507_),
    .Y(_1895_));
 sky130_fd_sc_hd__o31ai_2 _4245_ (.A1(_1870_),
    .A2(_1875_),
    .A3(_1895_),
    .B1(_1844_),
    .Y(_1896_));
 sky130_fd_sc_hd__nand2_1 _4246_ (.A(net2188),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .Y(_1897_));
 sky130_fd_sc_hd__xor2_1 _4247_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .B(_1896_),
    .X(_1898_));
 sky130_fd_sc_hd__and3b_1 _4248_ (.A_N(net2232),
    .B(net2354),
    .C(net2293),
    .X(_1899_));
 sky130_fd_sc_hd__inv_2 _4249_ (.A(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__nand2b_4 _4250_ (.A_N(net2188),
    .B(net2346),
    .Y(_1901_));
 sky130_fd_sc_hd__nand2b_4 _4251_ (.A_N(net2346),
    .B(net2188),
    .Y(_1902_));
 sky130_fd_sc_hd__or3_4 _4252_ (.A(net2293),
    .B(net2354),
    .C(net2232),
    .X(_1903_));
 sky130_fd_sc_hd__o22a_1 _4253_ (.A1(_1900_),
    .A2(_1901_),
    .B1(_1902_),
    .B2(_1903_),
    .X(_1904_));
 sky130_fd_sc_hd__or3b_4 _4254_ (.A(net2354),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .C_N(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .X(_1905_));
 sky130_fd_sc_hd__o21a_1 _4255_ (.A1(_1902_),
    .A2(_1905_),
    .B1(_1904_),
    .X(_1906_));
 sky130_fd_sc_hd__or2_1 _4256_ (.A(_1900_),
    .B(_1902_),
    .X(_1907_));
 sky130_fd_sc_hd__mux2_1 _4257_ (.A0(_1906_),
    .A1(_1907_),
    .S(_1844_),
    .X(_1908_));
 sky130_fd_sc_hd__o31ai_2 _4258_ (.A1(net2232),
    .A2(net2189),
    .A3(_1898_),
    .B1(_1908_),
    .Y(_1909_));
 sky130_fd_sc_hd__a21oi_4 _4259_ (.A1(net2154),
    .A2(_1909_),
    .B1(net2108),
    .Y(_1910_));
 sky130_fd_sc_hd__mux2_1 _4260_ (.A0(net2307),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[3] ),
    .S(net377),
    .X(_1911_));
 sky130_fd_sc_hd__nor2_1 _4261_ (.A(net2263),
    .B(_1911_),
    .Y(_1912_));
 sky130_fd_sc_hd__and2_1 _4262_ (.A(net2263),
    .B(_1911_),
    .X(_1913_));
 sky130_fd_sc_hd__or2_1 _4263_ (.A(net2264),
    .B(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__mux2_1 _4264_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[2] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[2] ),
    .S(net377),
    .X(_1915_));
 sky130_fd_sc_hd__and2_1 _4265_ (.A(net2333),
    .B(_1915_),
    .X(_1916_));
 sky130_fd_sc_hd__and3_1 _4266_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[1] ),
    .B(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ),
    .C(net2370),
    .X(_1917_));
 sky130_fd_sc_hd__a21oi_1 _4267_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ),
    .A2(net378),
    .B1(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[1] ),
    .Y(_1918_));
 sky130_fd_sc_hd__or2_1 _4268_ (.A(_1917_),
    .B(_1918_),
    .X(_1919_));
 sky130_fd_sc_hd__nand3_1 _4269_ (.A(net2150),
    .B(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ),
    .C(net378),
    .Y(_1920_));
 sky130_fd_sc_hd__nor2_1 _4270_ (.A(_1919_),
    .B(net2151),
    .Y(_1921_));
 sky130_fd_sc_hd__or2_2 _4271_ (.A(_1917_),
    .B(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__nor2_1 _4272_ (.A(net2333),
    .B(_1915_),
    .Y(_1923_));
 sky130_fd_sc_hd__or2_1 _4273_ (.A(_1916_),
    .B(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__and2b_1 _4274_ (.A_N(_1924_),
    .B(_1922_),
    .X(_1925_));
 sky130_fd_sc_hd__or2_1 _4275_ (.A(_1916_),
    .B(_1925_),
    .X(_1926_));
 sky130_fd_sc_hd__o21ba_1 _4276_ (.A1(_1916_),
    .A2(_1925_),
    .B1_N(_1914_),
    .X(_1927_));
 sky130_fd_sc_hd__xnor2_1 _4277_ (.A(net2265),
    .B(_1926_),
    .Y(_1928_));
 sky130_fd_sc_hd__mux2_1 _4278_ (.A0(_1928_),
    .A1(net2052),
    .S(net181),
    .X(_1929_));
 sky130_fd_sc_hd__and2b_1 _4279_ (.A_N(_1922_),
    .B(_1924_),
    .X(_1930_));
 sky130_fd_sc_hd__nor2_1 _4280_ (.A(_1925_),
    .B(_1930_),
    .Y(_1931_));
 sky130_fd_sc_hd__mux2_4 _4281_ (.A0(_1931_),
    .A1(net2131),
    .S(net183),
    .X(_1932_));
 sky130_fd_sc_hd__inv_2 _4282_ (.A(_1932_),
    .Y(_1933_));
 sky130_fd_sc_hd__nand2_1 _4283_ (.A(_1929_),
    .B(_1932_),
    .Y(_1934_));
 sky130_fd_sc_hd__mux2_1 _4284_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[4] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[4] ),
    .S(net377),
    .X(_1935_));
 sky130_fd_sc_hd__nor2_1 _4285_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ),
    .B(_1935_),
    .Y(_1936_));
 sky130_fd_sc_hd__and2_1 _4286_ (.A(net2295),
    .B(_1935_),
    .X(_1937_));
 sky130_fd_sc_hd__or2_1 _4287_ (.A(_1936_),
    .B(_1937_),
    .X(_1938_));
 sky130_fd_sc_hd__o21ba_1 _4288_ (.A1(_1913_),
    .A2(_1927_),
    .B1_N(_1938_),
    .X(_1939_));
 sky130_fd_sc_hd__or3b_1 _4289_ (.A(_1913_),
    .B(_1927_),
    .C_N(_1938_),
    .X(_1940_));
 sky130_fd_sc_hd__and2b_1 _4290_ (.A_N(_1939_),
    .B(net2308),
    .X(_1941_));
 sky130_fd_sc_hd__mux2_1 _4291_ (.A0(_1941_),
    .A1(net2013),
    .S(net181),
    .X(_1942_));
 sky130_fd_sc_hd__nand2b_2 _4292_ (.A_N(_1934_),
    .B(_1942_),
    .Y(_1943_));
 sky130_fd_sc_hd__mux2_1 _4293_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[5] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[5] ),
    .S(net377),
    .X(_1944_));
 sky130_fd_sc_hd__nor2_1 _4294_ (.A(net2191),
    .B(_1944_),
    .Y(_1945_));
 sky130_fd_sc_hd__and2_1 _4295_ (.A(net2191),
    .B(_1944_),
    .X(_1946_));
 sky130_fd_sc_hd__or2_1 _4296_ (.A(_1945_),
    .B(_1946_),
    .X(_1947_));
 sky130_fd_sc_hd__o21ba_1 _4297_ (.A1(_1937_),
    .A2(_1939_),
    .B1_N(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__or3b_1 _4298_ (.A(net2296),
    .B(_1939_),
    .C_N(_1947_),
    .X(_1949_));
 sky130_fd_sc_hd__and2b_1 _4299_ (.A_N(_1948_),
    .B(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__mux2_1 _4300_ (.A0(_1950_),
    .A1(net2005),
    .S(net178),
    .X(_1951_));
 sky130_fd_sc_hd__inv_2 _4301_ (.A(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__mux2_1 _4302_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[6] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ),
    .S(net377),
    .X(_1953_));
 sky130_fd_sc_hd__nor2_1 _4303_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ),
    .B(_1953_),
    .Y(_1954_));
 sky130_fd_sc_hd__and2_1 _4304_ (.A(net2177),
    .B(_1953_),
    .X(_1955_));
 sky130_fd_sc_hd__or2_1 _4305_ (.A(_1954_),
    .B(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__o21ba_1 _4306_ (.A1(_1946_),
    .A2(_1948_),
    .B1_N(_1956_),
    .X(_1957_));
 sky130_fd_sc_hd__or3b_1 _4307_ (.A(net2192),
    .B(_1948_),
    .C_N(_1956_),
    .X(_1958_));
 sky130_fd_sc_hd__and2b_1 _4308_ (.A_N(_1957_),
    .B(net2193),
    .X(_1959_));
 sky130_fd_sc_hd__mux2_1 _4309_ (.A0(_1959_),
    .A1(net1982),
    .S(net178),
    .X(_1960_));
 sky130_fd_sc_hd__inv_2 _4310_ (.A(_1960_),
    .Y(_1961_));
 sky130_fd_sc_hd__or3_1 _4311_ (.A(_1943_),
    .B(_1952_),
    .C(_1961_),
    .X(_1962_));
 sky130_fd_sc_hd__mux2_1 _4312_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[7] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[7] ),
    .S(net377),
    .X(_1963_));
 sky130_fd_sc_hd__nor2_1 _4313_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ),
    .B(_1963_),
    .Y(_1964_));
 sky130_fd_sc_hd__and2_1 _4314_ (.A(net2184),
    .B(_1963_),
    .X(_1965_));
 sky130_fd_sc_hd__or2_1 _4315_ (.A(_1964_),
    .B(_1965_),
    .X(_1966_));
 sky130_fd_sc_hd__o21ba_1 _4316_ (.A1(net2178),
    .A2(_1957_),
    .B1_N(_1966_),
    .X(_1967_));
 sky130_fd_sc_hd__or3b_1 _4317_ (.A(net2178),
    .B(_1957_),
    .C_N(_1966_),
    .X(_1968_));
 sky130_fd_sc_hd__and2b_1 _4318_ (.A_N(_1967_),
    .B(net2179),
    .X(_1969_));
 sky130_fd_sc_hd__mux2_1 _4319_ (.A0(_1969_),
    .A1(net1969),
    .S(net175),
    .X(_1970_));
 sky130_fd_sc_hd__nand2b_1 _4320_ (.A_N(_1962_),
    .B(_1970_),
    .Y(_1971_));
 sky130_fd_sc_hd__mux2_1 _4321_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[8] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[8] ),
    .S(net378),
    .X(_1972_));
 sky130_fd_sc_hd__nor2_1 _4322_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ),
    .B(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__and2_1 _4323_ (.A(net2301),
    .B(_1972_),
    .X(_1974_));
 sky130_fd_sc_hd__or2_1 _4324_ (.A(_1973_),
    .B(_1974_),
    .X(_1975_));
 sky130_fd_sc_hd__o21ba_1 _4325_ (.A1(net2185),
    .A2(_1967_),
    .B1_N(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__or3b_1 _4326_ (.A(net2185),
    .B(_1967_),
    .C_N(_1975_),
    .X(_1977_));
 sky130_fd_sc_hd__nand2b_1 _4327_ (.A_N(_1976_),
    .B(net2186),
    .Y(_1978_));
 sky130_fd_sc_hd__inv_2 _4328_ (.A(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__mux2_1 _4329_ (.A0(_1979_),
    .A1(net2033),
    .S(net176),
    .X(_1980_));
 sky130_fd_sc_hd__nand2b_2 _4330_ (.A_N(_1971_),
    .B(_1980_),
    .Y(_1981_));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[9] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ),
    .S(net377),
    .X(_1982_));
 sky130_fd_sc_hd__nor2_1 _4332_ (.A(net2274),
    .B(_1982_),
    .Y(_1983_));
 sky130_fd_sc_hd__and2_1 _4333_ (.A(net2274),
    .B(_1982_),
    .X(_1984_));
 sky130_fd_sc_hd__or2_1 _4334_ (.A(_1983_),
    .B(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__o21ba_1 _4335_ (.A1(_1974_),
    .A2(_1976_),
    .B1_N(_1985_),
    .X(_1986_));
 sky130_fd_sc_hd__or3b_1 _4336_ (.A(net2302),
    .B(_1976_),
    .C_N(_1985_),
    .X(_1987_));
 sky130_fd_sc_hd__and2b_1 _4337_ (.A_N(_1986_),
    .B(_1987_),
    .X(_1988_));
 sky130_fd_sc_hd__mux2_1 _4338_ (.A0(_1988_),
    .A1(net2001),
    .S(net178),
    .X(_1989_));
 sky130_fd_sc_hd__and2b_1 _4339_ (.A_N(_1981_),
    .B(_1989_),
    .X(_1990_));
 sky130_fd_sc_hd__mux2_1 _4340_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[10] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[10] ),
    .S(net378),
    .X(_1991_));
 sky130_fd_sc_hd__nor2_1 _4341_ (.A(net2270),
    .B(_1991_),
    .Y(_1992_));
 sky130_fd_sc_hd__and2_1 _4342_ (.A(net2270),
    .B(_1991_),
    .X(_1993_));
 sky130_fd_sc_hd__or2_1 _4343_ (.A(_1992_),
    .B(_1993_),
    .X(_1994_));
 sky130_fd_sc_hd__o21ba_1 _4344_ (.A1(_1984_),
    .A2(_1986_),
    .B1_N(_1994_),
    .X(_1995_));
 sky130_fd_sc_hd__or3b_1 _4345_ (.A(net2275),
    .B(_1986_),
    .C_N(_1994_),
    .X(_1996_));
 sky130_fd_sc_hd__and2b_1 _4346_ (.A_N(_1995_),
    .B(_1996_),
    .X(_1997_));
 sky130_fd_sc_hd__mux2_1 _4347_ (.A0(_1997_),
    .A1(net2038),
    .S(net176),
    .X(_1998_));
 sky130_fd_sc_hd__and2_1 _4348_ (.A(_1990_),
    .B(_1998_),
    .X(_1999_));
 sky130_fd_sc_hd__mux2_1 _4349_ (.A0(net2289),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ),
    .S(net377),
    .X(_2000_));
 sky130_fd_sc_hd__nor2_1 _4350_ (.A(net2369),
    .B(_2000_),
    .Y(_2001_));
 sky130_fd_sc_hd__and2_1 _4351_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ),
    .B(net2290),
    .X(_2002_));
 sky130_fd_sc_hd__or2_1 _4352_ (.A(_2001_),
    .B(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__o21ba_1 _4353_ (.A1(_1993_),
    .A2(_1995_),
    .B1_N(_2003_),
    .X(_2004_));
 sky130_fd_sc_hd__or3b_1 _4354_ (.A(net2271),
    .B(_1995_),
    .C_N(_2003_),
    .X(_2005_));
 sky130_fd_sc_hd__and2b_1 _4355_ (.A_N(_2004_),
    .B(_2005_),
    .X(_2006_));
 sky130_fd_sc_hd__mux2_1 _4356_ (.A0(_2006_),
    .A1(net1996),
    .S(net176),
    .X(_2007_));
 sky130_fd_sc_hd__nand2_1 _4357_ (.A(_1999_),
    .B(_2007_),
    .Y(_2008_));
 sky130_fd_sc_hd__mux2_1 _4358_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[12] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ),
    .S(net377),
    .X(_2009_));
 sky130_fd_sc_hd__nor2_1 _4359_ (.A(net2223),
    .B(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__and2_1 _4360_ (.A(net2223),
    .B(_2009_),
    .X(_2011_));
 sky130_fd_sc_hd__or2_1 _4361_ (.A(_2010_),
    .B(_2011_),
    .X(_2012_));
 sky130_fd_sc_hd__o21ba_1 _4362_ (.A1(net2360),
    .A2(_2004_),
    .B1_N(_2012_),
    .X(_2013_));
 sky130_fd_sc_hd__or3b_1 _4363_ (.A(net2291),
    .B(_2004_),
    .C_N(_2012_),
    .X(_2014_));
 sky130_fd_sc_hd__and2b_1 _4364_ (.A_N(_2013_),
    .B(_2014_),
    .X(_2015_));
 sky130_fd_sc_hd__mux2_2 _4365_ (.A0(_2015_),
    .A1(net1949),
    .S(net175),
    .X(_2016_));
 sky130_fd_sc_hd__mux2_1 _4366_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[13] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ),
    .S(net377),
    .X(_2017_));
 sky130_fd_sc_hd__nor2_1 _4367_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ),
    .B(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__and2_1 _4368_ (.A(net2286),
    .B(_2017_),
    .X(_2019_));
 sky130_fd_sc_hd__or2_1 _4369_ (.A(_2018_),
    .B(_2019_),
    .X(_2020_));
 sky130_fd_sc_hd__o21ba_1 _4370_ (.A1(net2224),
    .A2(_2013_),
    .B1_N(_2020_),
    .X(_2021_));
 sky130_fd_sc_hd__or3b_1 _4371_ (.A(net2224),
    .B(_2013_),
    .C_N(_2020_),
    .X(_2022_));
 sky130_fd_sc_hd__and2b_1 _4372_ (.A_N(_2021_),
    .B(net2225),
    .X(_2023_));
 sky130_fd_sc_hd__mux2_2 _4373_ (.A0(_2023_),
    .A1(net2048),
    .S(net178),
    .X(_2024_));
 sky130_fd_sc_hd__nand3b_4 _4374_ (.A_N(_2008_),
    .B(_2016_),
    .C(_2024_),
    .Y(_2025_));
 sky130_fd_sc_hd__mux2_1 _4375_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[14] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[14] ),
    .S(net377),
    .X(_2026_));
 sky130_fd_sc_hd__nor2_1 _4376_ (.A(net2241),
    .B(_2026_),
    .Y(_2027_));
 sky130_fd_sc_hd__and2_1 _4377_ (.A(net2241),
    .B(_2026_),
    .X(_2028_));
 sky130_fd_sc_hd__or2_1 _4378_ (.A(_2027_),
    .B(_2028_),
    .X(_2029_));
 sky130_fd_sc_hd__o21ba_1 _4379_ (.A1(net2287),
    .A2(_2021_),
    .B1_N(_2029_),
    .X(_2030_));
 sky130_fd_sc_hd__or3b_1 _4380_ (.A(net2287),
    .B(_2021_),
    .C_N(_2029_),
    .X(_2031_));
 sky130_fd_sc_hd__nand2b_1 _4381_ (.A_N(_2030_),
    .B(net2288),
    .Y(_2032_));
 sky130_fd_sc_hd__inv_2 _4382_ (.A(_2032_),
    .Y(_2033_));
 sky130_fd_sc_hd__mux2_1 _4383_ (.A0(_2033_),
    .A1(net2028),
    .S(net178),
    .X(_2034_));
 sky130_fd_sc_hd__and2b_1 _4384_ (.A_N(_2025_),
    .B(_2034_),
    .X(_2035_));
 sky130_fd_sc_hd__mux2_1 _4385_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[15] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[15] ),
    .S(net377),
    .X(_2036_));
 sky130_fd_sc_hd__nor2_1 _4386_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ),
    .B(_2036_),
    .Y(_2037_));
 sky130_fd_sc_hd__and2_1 _4387_ (.A(net2279),
    .B(_2036_),
    .X(_2038_));
 sky130_fd_sc_hd__or2_1 _4388_ (.A(_2037_),
    .B(_2038_),
    .X(_2039_));
 sky130_fd_sc_hd__o21ba_1 _4389_ (.A1(_2028_),
    .A2(_2030_),
    .B1_N(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__or3b_1 _4390_ (.A(net2242),
    .B(_2030_),
    .C_N(_2039_),
    .X(_2041_));
 sky130_fd_sc_hd__and2b_1 _4391_ (.A_N(_2040_),
    .B(net2243),
    .X(_2042_));
 sky130_fd_sc_hd__mux2_1 _4392_ (.A0(_2042_),
    .A1(net2017),
    .S(net179),
    .X(_2043_));
 sky130_fd_sc_hd__and2_1 _4393_ (.A(_2035_),
    .B(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__mux2_1 _4394_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[16] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ),
    .S(net377),
    .X(_2045_));
 sky130_fd_sc_hd__nor2_1 _4395_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ),
    .B(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__and2_1 _4396_ (.A(net2252),
    .B(_2045_),
    .X(_2047_));
 sky130_fd_sc_hd__or2_1 _4397_ (.A(_2046_),
    .B(_2047_),
    .X(_2048_));
 sky130_fd_sc_hd__o21ba_1 _4398_ (.A1(_2038_),
    .A2(_2040_),
    .B1_N(_2048_),
    .X(_2049_));
 sky130_fd_sc_hd__or3b_1 _4399_ (.A(net2280),
    .B(_2040_),
    .C_N(_2048_),
    .X(_2050_));
 sky130_fd_sc_hd__and2b_1 _4400_ (.A_N(_2049_),
    .B(_2050_),
    .X(_2051_));
 sky130_fd_sc_hd__mux2_1 _4401_ (.A0(_2051_),
    .A1(net2042),
    .S(net178),
    .X(_2052_));
 sky130_fd_sc_hd__mux2_1 _4402_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[17] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ),
    .S(net377),
    .X(_2053_));
 sky130_fd_sc_hd__nor2_1 _4403_ (.A(net2209),
    .B(_2053_),
    .Y(_2054_));
 sky130_fd_sc_hd__and2_1 _4404_ (.A(net2209),
    .B(_2053_),
    .X(_2055_));
 sky130_fd_sc_hd__or2_1 _4405_ (.A(_2054_),
    .B(_2055_),
    .X(_2056_));
 sky130_fd_sc_hd__o21ba_1 _4406_ (.A1(net2253),
    .A2(_2049_),
    .B1_N(_2056_),
    .X(_2057_));
 sky130_fd_sc_hd__or3b_1 _4407_ (.A(net2253),
    .B(_2049_),
    .C_N(_2056_),
    .X(_2058_));
 sky130_fd_sc_hd__nand2b_1 _4408_ (.A_N(_2057_),
    .B(net2254),
    .Y(_2059_));
 sky130_fd_sc_hd__inv_2 _4409_ (.A(_2059_),
    .Y(_2060_));
 sky130_fd_sc_hd__mux2_1 _4410_ (.A0(_2060_),
    .A1(net2079),
    .S(net179),
    .X(_2061_));
 sky130_fd_sc_hd__and3_4 _4411_ (.A(_2044_),
    .B(_2052_),
    .C(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__mux2_1 _4412_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[18] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[18] ),
    .S(net377),
    .X(_2063_));
 sky130_fd_sc_hd__nor2_1 _4413_ (.A(net2248),
    .B(_2063_),
    .Y(_2064_));
 sky130_fd_sc_hd__and2_1 _4414_ (.A(net2248),
    .B(_2063_),
    .X(_2065_));
 sky130_fd_sc_hd__or2_1 _4415_ (.A(_2064_),
    .B(_2065_),
    .X(_2066_));
 sky130_fd_sc_hd__o21ba_1 _4416_ (.A1(_2055_),
    .A2(_2057_),
    .B1_N(_2066_),
    .X(_2067_));
 sky130_fd_sc_hd__or3b_1 _4417_ (.A(net2210),
    .B(_2057_),
    .C_N(_2066_),
    .X(_2068_));
 sky130_fd_sc_hd__and2b_1 _4418_ (.A_N(_2067_),
    .B(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__mux2_1 _4419_ (.A0(_2069_),
    .A1(net2030),
    .S(net182),
    .X(_2070_));
 sky130_fd_sc_hd__and2_1 _4420_ (.A(_2062_),
    .B(_2070_),
    .X(_2071_));
 sky130_fd_sc_hd__mux2_1 _4421_ (.A0(net2277),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[19] ),
    .S(net2257),
    .X(_2072_));
 sky130_fd_sc_hd__nor2_1 _4422_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ),
    .B(_2072_),
    .Y(_2073_));
 sky130_fd_sc_hd__and2_1 _4423_ (.A(net2273),
    .B(net2278),
    .X(_2074_));
 sky130_fd_sc_hd__or2_1 _4424_ (.A(_2073_),
    .B(_2074_),
    .X(_2075_));
 sky130_fd_sc_hd__o21ba_1 _4425_ (.A1(_2065_),
    .A2(_2067_),
    .B1_N(_2075_),
    .X(_2076_));
 sky130_fd_sc_hd__or3b_1 _4426_ (.A(net2249),
    .B(_2067_),
    .C_N(_2075_),
    .X(_2077_));
 sky130_fd_sc_hd__and2b_1 _4427_ (.A_N(_2076_),
    .B(net2250),
    .X(_2078_));
 sky130_fd_sc_hd__mux2_2 _4428_ (.A0(_2078_),
    .A1(net1333),
    .S(net184),
    .X(_2079_));
 sky130_fd_sc_hd__nand2_1 _4429_ (.A(_2071_),
    .B(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__mux2_1 _4430_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[20] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[20] ),
    .S(net378),
    .X(_2081_));
 sky130_fd_sc_hd__nor2_1 _4431_ (.A(net2160),
    .B(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__and2_1 _4432_ (.A(net2160),
    .B(_2081_),
    .X(_2083_));
 sky130_fd_sc_hd__or2_4 _4433_ (.A(_2082_),
    .B(_2083_),
    .X(_2084_));
 sky130_fd_sc_hd__o21ba_4 _4434_ (.A1(_2074_),
    .A2(_2076_),
    .B1_N(_2084_),
    .X(_2085_));
 sky130_fd_sc_hd__or3b_1 _4435_ (.A(_2074_),
    .B(_2076_),
    .C_N(_2084_),
    .X(_2086_));
 sky130_fd_sc_hd__nand2b_2 _4436_ (.A_N(_2085_),
    .B(_2086_),
    .Y(_2087_));
 sky130_fd_sc_hd__inv_2 _4437_ (.A(_2087_),
    .Y(_2088_));
 sky130_fd_sc_hd__mux2_2 _4438_ (.A0(_2088_),
    .A1(net735),
    .S(net183),
    .X(_2089_));
 sky130_fd_sc_hd__and3_4 _4439_ (.A(_2071_),
    .B(_2079_),
    .C(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__mux2_1 _4440_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[21] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[21] ),
    .S(net378),
    .X(_2091_));
 sky130_fd_sc_hd__nor2_1 _4441_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ),
    .B(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__and2_1 _4442_ (.A(net2238),
    .B(_2091_),
    .X(_2093_));
 sky130_fd_sc_hd__or2_1 _4443_ (.A(_2092_),
    .B(_2093_),
    .X(_2094_));
 sky130_fd_sc_hd__o21ba_1 _4444_ (.A1(_2083_),
    .A2(_2085_),
    .B1_N(_2094_),
    .X(_2095_));
 sky130_fd_sc_hd__or3b_1 _4445_ (.A(net2161),
    .B(_2085_),
    .C_N(_2094_),
    .X(_2096_));
 sky130_fd_sc_hd__and2b_1 _4446_ (.A_N(_2095_),
    .B(net2162),
    .X(_2097_));
 sky130_fd_sc_hd__mux2_1 _4447_ (.A0(_2097_),
    .A1(net1828),
    .S(net174),
    .X(_2098_));
 sky130_fd_sc_hd__and2_4 _4448_ (.A(_2090_),
    .B(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__mux2_4 _4449_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[22] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ),
    .S(net377),
    .X(_2100_));
 sky130_fd_sc_hd__nor2_1 _4450_ (.A(net2200),
    .B(_2100_),
    .Y(_2101_));
 sky130_fd_sc_hd__and2_1 _4451_ (.A(net2200),
    .B(_2100_),
    .X(_2102_));
 sky130_fd_sc_hd__or2_1 _4452_ (.A(_2101_),
    .B(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__o21ba_1 _4453_ (.A1(net2239),
    .A2(_2095_),
    .B1_N(_2103_),
    .X(_2104_));
 sky130_fd_sc_hd__or3b_1 _4454_ (.A(net2239),
    .B(_2095_),
    .C_N(_2103_),
    .X(_2105_));
 sky130_fd_sc_hd__nand2b_1 _4455_ (.A_N(_2104_),
    .B(_2105_),
    .Y(_2106_));
 sky130_fd_sc_hd__inv_2 _4456_ (.A(_2106_),
    .Y(_2107_));
 sky130_fd_sc_hd__mux2_2 _4457_ (.A0(_2107_),
    .A1(net2016),
    .S(net173),
    .X(_2108_));
 sky130_fd_sc_hd__mux2_1 _4458_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[23] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[23] ),
    .S(net378),
    .X(_2109_));
 sky130_fd_sc_hd__nor2_1 _4459_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ),
    .B(_2109_),
    .Y(_2110_));
 sky130_fd_sc_hd__and2_1 _4460_ (.A(net2211),
    .B(_2109_),
    .X(_2111_));
 sky130_fd_sc_hd__or2_1 _4461_ (.A(_2110_),
    .B(_2111_),
    .X(_2112_));
 sky130_fd_sc_hd__o21ba_1 _4462_ (.A1(_2102_),
    .A2(_2104_),
    .B1_N(_2112_),
    .X(_2113_));
 sky130_fd_sc_hd__or3b_1 _4463_ (.A(_2102_),
    .B(_2104_),
    .C_N(_2112_),
    .X(_2114_));
 sky130_fd_sc_hd__and2b_1 _4464_ (.A_N(_2113_),
    .B(net2201),
    .X(_2115_));
 sky130_fd_sc_hd__mux2_1 _4465_ (.A0(_2115_),
    .A1(net661),
    .S(net173),
    .X(_2116_));
 sky130_fd_sc_hd__and3_1 _4466_ (.A(_2099_),
    .B(_2108_),
    .C(_2116_),
    .X(_2117_));
 sky130_fd_sc_hd__mux2_1 _4467_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[24] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ),
    .S(net378),
    .X(_2118_));
 sky130_fd_sc_hd__nor2_1 _4468_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ),
    .B(_2118_),
    .Y(_2119_));
 sky130_fd_sc_hd__and2_1 _4469_ (.A(net2123),
    .B(_2118_),
    .X(_2120_));
 sky130_fd_sc_hd__or2_1 _4470_ (.A(_2119_),
    .B(_2120_),
    .X(_2121_));
 sky130_fd_sc_hd__o21ba_1 _4471_ (.A1(_2111_),
    .A2(_2113_),
    .B1_N(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__or3b_1 _4472_ (.A(net2212),
    .B(_2113_),
    .C_N(_2121_),
    .X(_2123_));
 sky130_fd_sc_hd__and2b_1 _4473_ (.A_N(_2122_),
    .B(net2213),
    .X(_2124_));
 sky130_fd_sc_hd__mux2_1 _4474_ (.A0(_2124_),
    .A1(net2072),
    .S(net177),
    .X(_2125_));
 sky130_fd_sc_hd__and2_1 _4475_ (.A(_2117_),
    .B(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__mux2_1 _4476_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[25] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[25] ),
    .S(net378),
    .X(_2127_));
 sky130_fd_sc_hd__nor2_1 _4477_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ),
    .B(_2127_),
    .Y(_2128_));
 sky130_fd_sc_hd__and2_1 _4478_ (.A(net2216),
    .B(_2127_),
    .X(_2129_));
 sky130_fd_sc_hd__or2_1 _4479_ (.A(_2128_),
    .B(_2129_),
    .X(_2130_));
 sky130_fd_sc_hd__o21ba_1 _4480_ (.A1(net2124),
    .A2(_2122_),
    .B1_N(_2130_),
    .X(_2131_));
 sky130_fd_sc_hd__or3b_1 _4481_ (.A(net2124),
    .B(_2122_),
    .C_N(_2130_),
    .X(_2132_));
 sky130_fd_sc_hd__and2b_1 _4482_ (.A_N(_2131_),
    .B(net2125),
    .X(_2133_));
 sky130_fd_sc_hd__mux2_1 _4483_ (.A0(_2133_),
    .A1(net2098),
    .S(net172),
    .X(_2134_));
 sky130_fd_sc_hd__and3_1 _4484_ (.A(_2117_),
    .B(_2125_),
    .C(_2134_),
    .X(_2135_));
 sky130_fd_sc_hd__mux2_1 _4485_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[26] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[26] ),
    .S(net378),
    .X(_2136_));
 sky130_fd_sc_hd__nor2_1 _4486_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ),
    .B(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__and2_1 _4487_ (.A(net2305),
    .B(_2136_),
    .X(_2138_));
 sky130_fd_sc_hd__or2_1 _4488_ (.A(_2137_),
    .B(_2138_),
    .X(_2139_));
 sky130_fd_sc_hd__o21ba_1 _4489_ (.A1(_2129_),
    .A2(_2131_),
    .B1_N(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__or3b_1 _4490_ (.A(net2217),
    .B(_2131_),
    .C_N(_2139_),
    .X(_2141_));
 sky130_fd_sc_hd__and2b_1 _4491_ (.A_N(_2140_),
    .B(net2218),
    .X(_2142_));
 sky130_fd_sc_hd__mux2_1 _4492_ (.A0(_2142_),
    .A1(net2087),
    .S(net172),
    .X(_2143_));
 sky130_fd_sc_hd__and2_1 _4493_ (.A(_2135_),
    .B(_2143_),
    .X(_2144_));
 sky130_fd_sc_hd__mux2_1 _4494_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[27] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[27] ),
    .S(net378),
    .X(_2145_));
 sky130_fd_sc_hd__nor2_1 _4495_ (.A(net2282),
    .B(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__and2_1 _4496_ (.A(net2282),
    .B(_2145_),
    .X(_2147_));
 sky130_fd_sc_hd__or2_1 _4497_ (.A(_2146_),
    .B(_2147_),
    .X(_2148_));
 sky130_fd_sc_hd__o21ba_1 _4498_ (.A1(_2138_),
    .A2(_2140_),
    .B1_N(_2148_),
    .X(_2149_));
 sky130_fd_sc_hd__or3b_1 _4499_ (.A(net2306),
    .B(_2140_),
    .C_N(_2148_),
    .X(_2150_));
 sky130_fd_sc_hd__and2b_1 _4500_ (.A_N(_2149_),
    .B(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__mux2_1 _4501_ (.A0(_2151_),
    .A1(net2060),
    .S(net173),
    .X(_2152_));
 sky130_fd_sc_hd__and3_2 _4502_ (.A(_2135_),
    .B(_2143_),
    .C(_2152_),
    .X(_2153_));
 sky130_fd_sc_hd__mux2_1 _4503_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[28] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[28] ),
    .S(net378),
    .X(_2154_));
 sky130_fd_sc_hd__nor2_1 _4504_ (.A(net2227),
    .B(_2154_),
    .Y(_2155_));
 sky130_fd_sc_hd__and2_1 _4505_ (.A(net2227),
    .B(_2154_),
    .X(_2156_));
 sky130_fd_sc_hd__or2_1 _4506_ (.A(_2155_),
    .B(_2156_),
    .X(_2157_));
 sky130_fd_sc_hd__o21ba_1 _4507_ (.A1(_2147_),
    .A2(_2149_),
    .B1_N(_2157_),
    .X(_2158_));
 sky130_fd_sc_hd__or3b_1 _4508_ (.A(net2283),
    .B(_2149_),
    .C_N(_2157_),
    .X(_2159_));
 sky130_fd_sc_hd__and2b_1 _4509_ (.A_N(_2158_),
    .B(net2284),
    .X(_2160_));
 sky130_fd_sc_hd__mux2_1 _4510_ (.A0(_2160_),
    .A1(net2043),
    .S(net171),
    .X(_2161_));
 sky130_fd_sc_hd__and2_1 _4511_ (.A(_2153_),
    .B(_2161_),
    .X(_2162_));
 sky130_fd_sc_hd__mux2_1 _4512_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[29] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[29] ),
    .S(net378),
    .X(_2163_));
 sky130_fd_sc_hd__nor2_1 _4513_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ),
    .B(_2163_),
    .Y(_2164_));
 sky130_fd_sc_hd__and2_1 _4514_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ),
    .B(_2163_),
    .X(_2165_));
 sky130_fd_sc_hd__or2_1 _4515_ (.A(_2164_),
    .B(_2165_),
    .X(_2166_));
 sky130_fd_sc_hd__o21ba_1 _4516_ (.A1(_2156_),
    .A2(_2158_),
    .B1_N(_2166_),
    .X(_2167_));
 sky130_fd_sc_hd__or3b_1 _4517_ (.A(net2228),
    .B(_2158_),
    .C_N(_2166_),
    .X(_2168_));
 sky130_fd_sc_hd__and2b_1 _4518_ (.A_N(_2167_),
    .B(net2229),
    .X(_2169_));
 sky130_fd_sc_hd__mux2_1 _4519_ (.A0(_2169_),
    .A1(net2049),
    .S(net171),
    .X(_2170_));
 sky130_fd_sc_hd__and3_1 _4520_ (.A(_2153_),
    .B(_2161_),
    .C(_2170_),
    .X(_2171_));
 sky130_fd_sc_hd__mux2_1 _4521_ (.A0(\U_DATAPATH.U_ID_EX.o_pc_EX[30] ),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ),
    .S(net378),
    .X(_2172_));
 sky130_fd_sc_hd__xnor2_1 _4522_ (.A(net2259),
    .B(_2172_),
    .Y(_2173_));
 sky130_fd_sc_hd__o21ba_1 _4523_ (.A1(_2165_),
    .A2(_2167_),
    .B1_N(net2260),
    .X(_2174_));
 sky130_fd_sc_hd__or3b_1 _4524_ (.A(_2165_),
    .B(_2167_),
    .C_N(net2260),
    .X(_2175_));
 sky130_fd_sc_hd__and2b_1 _4525_ (.A_N(_2174_),
    .B(net2261),
    .X(_2176_));
 sky130_fd_sc_hd__mux2_1 _4526_ (.A0(_2176_),
    .A1(net2070),
    .S(net174),
    .X(_2177_));
 sky130_fd_sc_hd__and2_4 _4527_ (.A(_2171_),
    .B(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__a21o_1 _4528_ (.A1(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ),
    .A2(_2172_),
    .B1(_2174_),
    .X(_2179_));
 sky130_fd_sc_hd__xnor2_2 _4529_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ),
    .B(_2179_),
    .Y(_2180_));
 sky130_fd_sc_hd__mux2_1 _4530_ (.A0(net2022),
    .A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ),
    .S(net378),
    .X(_2181_));
 sky130_fd_sc_hd__xnor2_1 _4531_ (.A(_2180_),
    .B(net2023),
    .Y(_2182_));
 sky130_fd_sc_hd__mux2_1 _4532_ (.A0(net2024),
    .A1(net1850),
    .S(net173),
    .X(_2183_));
 sky130_fd_sc_hd__or2_1 _4533_ (.A(net394),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .X(_2184_));
 sky130_fd_sc_hd__nand2_1 _4534_ (.A(net394),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .Y(_2185_));
 sky130_fd_sc_hd__or2_1 _4535_ (.A(net404),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .X(_2186_));
 sky130_fd_sc_hd__nand2_1 _4536_ (.A(net404),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .Y(_2187_));
 sky130_fd_sc_hd__a22o_1 _4537_ (.A1(_2184_),
    .A2(_2185_),
    .B1(_2186_),
    .B2(_2187_),
    .X(_2188_));
 sky130_fd_sc_hd__or2_1 _4538_ (.A(net382),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .X(_2189_));
 sky130_fd_sc_hd__nand2_1 _4539_ (.A(net382),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .Y(_2190_));
 sky130_fd_sc_hd__or2_1 _4540_ (.A(net387),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .X(_2191_));
 sky130_fd_sc_hd__nand2_1 _4541_ (.A(net387),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .Y(_2192_));
 sky130_fd_sc_hd__a22o_1 _4542_ (.A1(_2189_),
    .A2(_2190_),
    .B1(_2191_),
    .B2(_2192_),
    .X(_2193_));
 sky130_fd_sc_hd__or2_1 _4543_ (.A(net433),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .X(_2194_));
 sky130_fd_sc_hd__nand2_1 _4544_ (.A(net433),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .Y(_2195_));
 sky130_fd_sc_hd__or2_1 _4545_ (.A(net409),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .X(_2196_));
 sky130_fd_sc_hd__nand2_1 _4546_ (.A(net409),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .Y(_2197_));
 sky130_fd_sc_hd__or2_1 _4547_ (.A(net425),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .X(_2198_));
 sky130_fd_sc_hd__nand2_1 _4548_ (.A(net425),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .Y(_2199_));
 sky130_fd_sc_hd__or2_1 _4549_ (.A(net414),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .X(_2200_));
 sky130_fd_sc_hd__nand2_1 _4550_ (.A(net414),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .Y(_2201_));
 sky130_fd_sc_hd__a22o_1 _4551_ (.A1(_2194_),
    .A2(_2195_),
    .B1(_2198_),
    .B2(_2199_),
    .X(_2202_));
 sky130_fd_sc_hd__a22o_1 _4552_ (.A1(_2196_),
    .A2(_2197_),
    .B1(_2200_),
    .B2(_2201_),
    .X(_2203_));
 sky130_fd_sc_hd__o22a_4 _4553_ (.A1(_2188_),
    .A2(_2193_),
    .B1(_2202_),
    .B2(_2203_),
    .X(_2204_));
 sky130_fd_sc_hd__nor3b_4 _4554_ (.A(net1435),
    .B(_2204_),
    .C_N(net2031),
    .Y(_2205_));
 sky130_fd_sc_hd__or3b_2 _4555_ (.A(net1435),
    .B(_2204_),
    .C_N(net2031),
    .X(_2206_));
 sky130_fd_sc_hd__nor2_1 _4556_ (.A(_2178_),
    .B(net295),
    .Y(_2207_));
 sky130_fd_sc_hd__nand2_1 _4557_ (.A(_2178_),
    .B(_2183_),
    .Y(_2208_));
 sky130_fd_sc_hd__o21a_1 _4558_ (.A1(_2178_),
    .A2(_2183_),
    .B1(net280),
    .X(_2209_));
 sky130_fd_sc_hd__a22o_1 _4559_ (.A1(net1850),
    .A2(net294),
    .B1(_2208_),
    .B2(_2209_),
    .X(_1273_));
 sky130_fd_sc_hd__or2_1 _4560_ (.A(_2171_),
    .B(_2177_),
    .X(_2210_));
 sky130_fd_sc_hd__a22o_1 _4561_ (.A1(net2070),
    .A2(net295),
    .B1(_2207_),
    .B2(_2210_),
    .X(_1272_));
 sky130_fd_sc_hd__or2_1 _4562_ (.A(_2162_),
    .B(_2170_),
    .X(_2211_));
 sky130_fd_sc_hd__nor2_1 _4563_ (.A(_2171_),
    .B(net295),
    .Y(_2212_));
 sky130_fd_sc_hd__a22o_1 _4564_ (.A1(net2049),
    .A2(net295),
    .B1(_2211_),
    .B2(_2212_),
    .X(_1271_));
 sky130_fd_sc_hd__or2_1 _4565_ (.A(_2153_),
    .B(_2161_),
    .X(_2213_));
 sky130_fd_sc_hd__nor2_1 _4566_ (.A(_2162_),
    .B(net295),
    .Y(_2214_));
 sky130_fd_sc_hd__a22o_1 _4567_ (.A1(net2043),
    .A2(net295),
    .B1(_2213_),
    .B2(_2214_),
    .X(_1270_));
 sky130_fd_sc_hd__or2_1 _4568_ (.A(_2144_),
    .B(_2152_),
    .X(_2215_));
 sky130_fd_sc_hd__nor2_1 _4569_ (.A(_2153_),
    .B(net293),
    .Y(_2216_));
 sky130_fd_sc_hd__a22o_1 _4570_ (.A1(net2060),
    .A2(net293),
    .B1(_2215_),
    .B2(_2216_),
    .X(_1269_));
 sky130_fd_sc_hd__or2_1 _4571_ (.A(_2135_),
    .B(_2143_),
    .X(_2217_));
 sky130_fd_sc_hd__nor2_1 _4572_ (.A(_2144_),
    .B(net293),
    .Y(_2218_));
 sky130_fd_sc_hd__a22o_1 _4573_ (.A1(net2087),
    .A2(net293),
    .B1(_2217_),
    .B2(_2218_),
    .X(_1268_));
 sky130_fd_sc_hd__or2_1 _4574_ (.A(_2126_),
    .B(_2134_),
    .X(_2219_));
 sky130_fd_sc_hd__nor2_1 _4575_ (.A(_2135_),
    .B(net294),
    .Y(_2220_));
 sky130_fd_sc_hd__a22o_1 _4576_ (.A1(net2098),
    .A2(net293),
    .B1(_2219_),
    .B2(_2220_),
    .X(_1267_));
 sky130_fd_sc_hd__or2_1 _4577_ (.A(_2117_),
    .B(_2125_),
    .X(_2221_));
 sky130_fd_sc_hd__nor2_1 _4578_ (.A(_2126_),
    .B(net293),
    .Y(_2222_));
 sky130_fd_sc_hd__a22o_1 _4579_ (.A1(net2072),
    .A2(net293),
    .B1(_2221_),
    .B2(_2222_),
    .X(_1266_));
 sky130_fd_sc_hd__a31o_1 _4580_ (.A1(_2090_),
    .A2(_2098_),
    .A3(_2108_),
    .B1(_2116_),
    .X(_2223_));
 sky130_fd_sc_hd__nor2_1 _4581_ (.A(_2117_),
    .B(net294),
    .Y(_2224_));
 sky130_fd_sc_hd__a22o_1 _4582_ (.A1(net661),
    .A2(net294),
    .B1(_2223_),
    .B2(_2224_),
    .X(_1265_));
 sky130_fd_sc_hd__or2_1 _4583_ (.A(_2099_),
    .B(_2108_),
    .X(_2225_));
 sky130_fd_sc_hd__a21oi_1 _4584_ (.A1(_2099_),
    .A2(_2108_),
    .B1(net294),
    .Y(_2226_));
 sky130_fd_sc_hd__a22o_1 _4585_ (.A1(net2016),
    .A2(net294),
    .B1(_2225_),
    .B2(_2226_),
    .X(_1264_));
 sky130_fd_sc_hd__or2_1 _4586_ (.A(_2090_),
    .B(_2098_),
    .X(_2227_));
 sky130_fd_sc_hd__nor2_1 _4587_ (.A(_2099_),
    .B(net294),
    .Y(_2228_));
 sky130_fd_sc_hd__a22o_1 _4588_ (.A1(net1828),
    .A2(net294),
    .B1(_2227_),
    .B2(_2228_),
    .X(_1263_));
 sky130_fd_sc_hd__a31o_1 _4589_ (.A1(_2062_),
    .A2(_2070_),
    .A3(_2079_),
    .B1(_2089_),
    .X(_2229_));
 sky130_fd_sc_hd__nor2_1 _4590_ (.A(_2090_),
    .B(net302),
    .Y(_2230_));
 sky130_fd_sc_hd__a22o_1 _4591_ (.A1(net735),
    .A2(net301),
    .B1(_2229_),
    .B2(_2230_),
    .X(_1262_));
 sky130_fd_sc_hd__and2_1 _4592_ (.A(net1333),
    .B(net301),
    .X(_2231_));
 sky130_fd_sc_hd__or2_1 _4593_ (.A(_2071_),
    .B(_2079_),
    .X(_2232_));
 sky130_fd_sc_hd__a31o_1 _4594_ (.A1(_2080_),
    .A2(net289),
    .A3(_2232_),
    .B1(_2231_),
    .X(_1261_));
 sky130_fd_sc_hd__or2_1 _4595_ (.A(_2062_),
    .B(_2070_),
    .X(_2233_));
 sky130_fd_sc_hd__nor2_1 _4596_ (.A(_2071_),
    .B(net301),
    .Y(_2234_));
 sky130_fd_sc_hd__a22o_1 _4597_ (.A1(net2030),
    .A2(net302),
    .B1(_2233_),
    .B2(_2234_),
    .X(_1260_));
 sky130_fd_sc_hd__a21oi_1 _4598_ (.A1(_2044_),
    .A2(_2052_),
    .B1(_2061_),
    .Y(_2235_));
 sky130_fd_sc_hd__nor2_1 _4599_ (.A(_2062_),
    .B(_2235_),
    .Y(_2236_));
 sky130_fd_sc_hd__mux2_1 _4600_ (.A0(net2079),
    .A1(_2236_),
    .S(net285),
    .X(_1259_));
 sky130_fd_sc_hd__xor2_1 _4601_ (.A(_2044_),
    .B(_2052_),
    .X(_2237_));
 sky130_fd_sc_hd__mux2_1 _4602_ (.A0(net2042),
    .A1(_2237_),
    .S(net285),
    .X(_1258_));
 sky130_fd_sc_hd__or2_1 _4603_ (.A(_2035_),
    .B(_2043_),
    .X(_2238_));
 sky130_fd_sc_hd__nor2_1 _4604_ (.A(_2044_),
    .B(net300),
    .Y(_2239_));
 sky130_fd_sc_hd__a22o_1 _4605_ (.A1(net2017),
    .A2(net300),
    .B1(_2238_),
    .B2(_2239_),
    .X(_1257_));
 sky130_fd_sc_hd__nand2b_1 _4606_ (.A_N(_2034_),
    .B(_2025_),
    .Y(_2240_));
 sky130_fd_sc_hd__nor2_1 _4607_ (.A(_2035_),
    .B(net299),
    .Y(_2241_));
 sky130_fd_sc_hd__a22o_1 _4608_ (.A1(net2028),
    .A2(net299),
    .B1(_2240_),
    .B2(_2241_),
    .X(_1256_));
 sky130_fd_sc_hd__and2_1 _4609_ (.A(net2048),
    .B(net297),
    .X(_2242_));
 sky130_fd_sc_hd__a31o_1 _4610_ (.A1(_1999_),
    .A2(_2007_),
    .A3(_2016_),
    .B1(_2024_),
    .X(_2243_));
 sky130_fd_sc_hd__a31o_1 _4611_ (.A1(_2025_),
    .A2(net277),
    .A3(_2243_),
    .B1(_2242_),
    .X(_1255_));
 sky130_fd_sc_hd__xnor2_1 _4612_ (.A(_2008_),
    .B(_2016_),
    .Y(_2244_));
 sky130_fd_sc_hd__mux2_1 _4613_ (.A0(net1949),
    .A1(_2244_),
    .S(net278),
    .X(_1254_));
 sky130_fd_sc_hd__and2_1 _4614_ (.A(net1996),
    .B(net296),
    .X(_2245_));
 sky130_fd_sc_hd__or2_1 _4615_ (.A(_1999_),
    .B(_2007_),
    .X(_2246_));
 sky130_fd_sc_hd__a31o_1 _4616_ (.A1(_2008_),
    .A2(net277),
    .A3(_2246_),
    .B1(_2245_),
    .X(_1253_));
 sky130_fd_sc_hd__or2_1 _4617_ (.A(_1990_),
    .B(_1998_),
    .X(_2247_));
 sky130_fd_sc_hd__nor2_1 _4618_ (.A(_1999_),
    .B(net296),
    .Y(_2248_));
 sky130_fd_sc_hd__a22o_1 _4619_ (.A1(net2038),
    .A2(net296),
    .B1(_2247_),
    .B2(_2248_),
    .X(_1252_));
 sky130_fd_sc_hd__xnor2_1 _4620_ (.A(_1981_),
    .B(_1989_),
    .Y(_2249_));
 sky130_fd_sc_hd__mux2_1 _4621_ (.A0(net2001),
    .A1(_2249_),
    .S(net282),
    .X(_1251_));
 sky130_fd_sc_hd__and2_1 _4622_ (.A(net2033),
    .B(net297),
    .X(_2250_));
 sky130_fd_sc_hd__nand2b_1 _4623_ (.A_N(_1980_),
    .B(_1971_),
    .Y(_2251_));
 sky130_fd_sc_hd__a31o_1 _4624_ (.A1(_1981_),
    .A2(net282),
    .A3(_2251_),
    .B1(_2250_),
    .X(_1250_));
 sky130_fd_sc_hd__and2_1 _4625_ (.A(net1969),
    .B(net296),
    .X(_2252_));
 sky130_fd_sc_hd__nand2b_1 _4626_ (.A_N(_1970_),
    .B(_1962_),
    .Y(_2253_));
 sky130_fd_sc_hd__a31o_1 _4627_ (.A1(_1971_),
    .A2(net278),
    .A3(_2253_),
    .B1(_2252_),
    .X(_1249_));
 sky130_fd_sc_hd__and2_1 _4628_ (.A(net1982),
    .B(net299),
    .X(_2254_));
 sky130_fd_sc_hd__o21ai_1 _4629_ (.A1(net2014),
    .A2(_1952_),
    .B1(_1961_),
    .Y(_2255_));
 sky130_fd_sc_hd__a31o_1 _4630_ (.A1(_1962_),
    .A2(net282),
    .A3(_2255_),
    .B1(_2254_),
    .X(_1248_));
 sky130_fd_sc_hd__xnor2_1 _4631_ (.A(_1943_),
    .B(_1951_),
    .Y(_2256_));
 sky130_fd_sc_hd__mux2_1 _4632_ (.A0(net2005),
    .A1(net2015),
    .S(net282),
    .X(_1247_));
 sky130_fd_sc_hd__and2_1 _4633_ (.A(net2013),
    .B(net301),
    .X(_2257_));
 sky130_fd_sc_hd__a21o_1 _4634_ (.A1(_1929_),
    .A2(_1932_),
    .B1(_1942_),
    .X(_2258_));
 sky130_fd_sc_hd__a31o_1 _4635_ (.A1(net2014),
    .A2(net288),
    .A3(_2258_),
    .B1(_2257_),
    .X(_1246_));
 sky130_fd_sc_hd__and2_1 _4636_ (.A(net2052),
    .B(net301),
    .X(_2259_));
 sky130_fd_sc_hd__or2_1 _4637_ (.A(_1929_),
    .B(_1932_),
    .X(_2260_));
 sky130_fd_sc_hd__a31o_1 _4638_ (.A1(_1934_),
    .A2(net288),
    .A3(_2260_),
    .B1(_2259_),
    .X(_1245_));
 sky130_fd_sc_hd__mux2_1 _4639_ (.A0(net2131),
    .A1(_1933_),
    .S(net289),
    .X(_1244_));
 sky130_fd_sc_hd__and2_1 _4640_ (.A(\U_DATAPATH.U_EX_MEM.o_mem_write_M ),
    .B(net449),
    .X(_1016_));
 sky130_fd_sc_hd__and2_1 _4641_ (.A(net444),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[31] ),
    .X(_1015_));
 sky130_fd_sc_hd__and2_1 _4642_ (.A(net462),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[30] ),
    .X(_1014_));
 sky130_fd_sc_hd__and2_1 _4643_ (.A(net439),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[29] ),
    .X(_1013_));
 sky130_fd_sc_hd__and2_1 _4644_ (.A(net441),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[28] ),
    .X(_1012_));
 sky130_fd_sc_hd__and2_1 _4645_ (.A(net468),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[27] ),
    .X(_1011_));
 sky130_fd_sc_hd__and2_1 _4646_ (.A(net441),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[26] ),
    .X(_1010_));
 sky130_fd_sc_hd__and2_1 _4647_ (.A(net450),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[25] ),
    .X(_1009_));
 sky130_fd_sc_hd__and2_1 _4648_ (.A(net470),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[24] ),
    .X(_1008_));
 sky130_fd_sc_hd__and2_1 _4649_ (.A(net443),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[23] ),
    .X(_1007_));
 sky130_fd_sc_hd__and2_1 _4650_ (.A(net466),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[22] ),
    .X(_1006_));
 sky130_fd_sc_hd__and2_1 _4651_ (.A(net440),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[21] ),
    .X(_1005_));
 sky130_fd_sc_hd__and2_1 _4652_ (.A(net441),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[20] ),
    .X(_1004_));
 sky130_fd_sc_hd__and2_1 _4653_ (.A(net455),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[19] ),
    .X(_1003_));
 sky130_fd_sc_hd__and2_1 _4654_ (.A(net465),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[18] ),
    .X(_1002_));
 sky130_fd_sc_hd__and2_1 _4655_ (.A(net455),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[17] ),
    .X(_1001_));
 sky130_fd_sc_hd__and2_1 _4656_ (.A(net456),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[16] ),
    .X(_1000_));
 sky130_fd_sc_hd__and2_1 _4657_ (.A(net457),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[15] ),
    .X(_0999_));
 sky130_fd_sc_hd__and2_1 _4658_ (.A(net455),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[14] ),
    .X(_0998_));
 sky130_fd_sc_hd__and2_1 _4659_ (.A(net444),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[13] ),
    .X(_0997_));
 sky130_fd_sc_hd__and2_1 _4660_ (.A(net455),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[12] ),
    .X(_0996_));
 sky130_fd_sc_hd__and2_1 _4661_ (.A(net440),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[11] ),
    .X(_0995_));
 sky130_fd_sc_hd__and2_1 _4662_ (.A(net470),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[10] ),
    .X(_0994_));
 sky130_fd_sc_hd__and2_1 _4663_ (.A(net457),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[9] ),
    .X(_0993_));
 sky130_fd_sc_hd__and2_1 _4664_ (.A(net441),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[8] ),
    .X(_0992_));
 sky130_fd_sc_hd__and2_1 _4665_ (.A(net472),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[7] ),
    .X(_0991_));
 sky130_fd_sc_hd__and2_1 _4666_ (.A(net455),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[6] ),
    .X(_0990_));
 sky130_fd_sc_hd__and2_1 _4667_ (.A(net464),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[5] ),
    .X(_0989_));
 sky130_fd_sc_hd__and2_1 _4668_ (.A(net469),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[4] ),
    .X(_0988_));
 sky130_fd_sc_hd__and2_1 _4669_ (.A(net469),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[3] ),
    .X(_0987_));
 sky130_fd_sc_hd__and2_1 _4670_ (.A(net447),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[2] ),
    .X(_0986_));
 sky130_fd_sc_hd__and2_1 _4671_ (.A(net447),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[1] ),
    .X(_0985_));
 sky130_fd_sc_hd__and2_1 _4672_ (.A(net445),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[0] ),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _4673_ (.A0(net2078),
    .A1(_2183_),
    .S(net280),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _4674_ (.A0(net2082),
    .A1(_2177_),
    .S(net273),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _4675_ (.A0(net2097),
    .A1(_2170_),
    .S(net272),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _4676_ (.A0(net2076),
    .A1(_2161_),
    .S(net272),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _4677_ (.A0(net2095),
    .A1(_2152_),
    .S(net276),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _4678_ (.A0(net2102),
    .A1(_2143_),
    .S(net275),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _4679_ (.A0(net2075),
    .A1(_2134_),
    .S(net275),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _4680_ (.A0(net2088),
    .A1(_2125_),
    .S(net280),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _4681_ (.A0(net2064),
    .A1(_2116_),
    .S(net275),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _4682_ (.A0(net2083),
    .A1(_2108_),
    .S(net281),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _4683_ (.A0(net2090),
    .A1(_2098_),
    .S(net276),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _4684_ (.A0(net2080),
    .A1(_2089_),
    .S(net291),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _4685_ (.A0(net2116),
    .A1(_2079_),
    .S(net286),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _4686_ (.A0(net2051),
    .A1(_2070_),
    .S(net289),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _4687_ (.A0(net2096),
    .A1(_2061_),
    .S(net285),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _4688_ (.A0(net2069),
    .A1(_2052_),
    .S(net283),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _4689_ (.A0(net2068),
    .A1(_2043_),
    .S(net285),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _4690_ (.A0(net2104),
    .A1(_2034_),
    .S(net285),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _4691_ (.A0(net2071),
    .A1(_2024_),
    .S(net283),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _4692_ (.A0(net2081),
    .A1(_2016_),
    .S(net278),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _4693_ (.A0(net2077),
    .A1(_2007_),
    .S(net277),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _4694_ (.A0(net2089),
    .A1(_1998_),
    .S(net279),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _4695_ (.A0(net2036),
    .A1(_1989_),
    .S(net283),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _4696_ (.A0(net2041),
    .A1(net2034),
    .S(net278),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _4697_ (.A0(net2063),
    .A1(_1970_),
    .S(net277),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _4698_ (.A0(net2026),
    .A1(_1960_),
    .S(net277),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _4699_ (.A0(net2053),
    .A1(_1951_),
    .S(net282),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _4700_ (.A0(net2037),
    .A1(_1942_),
    .S(net288),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _4701_ (.A0(net2117),
    .A1(_1929_),
    .S(net288),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _4702_ (.A0(net2099),
    .A1(_1932_),
    .S(net289),
    .X(_0292_));
 sky130_fd_sc_hd__nand2b_1 _4703_ (.A_N(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .B(net2197),
    .Y(_2261_));
 sky130_fd_sc_hd__nor3_1 _4704_ (.A(_1407_),
    .B(_1408_),
    .C(net2198),
    .Y(_2262_));
 sky130_fd_sc_hd__or3_2 _4705_ (.A(_1407_),
    .B(_1408_),
    .C(net2198),
    .X(_2263_));
 sky130_fd_sc_hd__and4bb_4 _4706_ (.A_N(net2234),
    .B_N(net2058),
    .C(net2073),
    .D(net2203),
    .X(_2264_));
 sky130_fd_sc_hd__or4b_2 _4707_ (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .B(net2058),
    .C(_1408_),
    .D_N(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .X(_2265_));
 sky130_fd_sc_hd__o21a_2 _4708_ (.A1(net2197),
    .A2(net2059),
    .B1(_2263_),
    .X(_2266_));
 sky130_fd_sc_hd__or2_4 _4709_ (.A(net2058),
    .B(net2073),
    .X(_2267_));
 sky130_fd_sc_hd__o31a_1 _4710_ (.A1(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .A2(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .A3(_2267_),
    .B1(_2266_),
    .X(_3744_));
 sky130_fd_sc_hd__mux4_1 _4711_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ),
    .S0(net405),
    .S1(net395),
    .X(_2268_));
 sky130_fd_sc_hd__mux4_1 _4712_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ),
    .S0(net405),
    .S1(net395),
    .X(_2269_));
 sky130_fd_sc_hd__mux2_1 _4713_ (.A0(_2268_),
    .A1(_2269_),
    .S(net386),
    .X(_2270_));
 sky130_fd_sc_hd__mux4_1 _4714_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ),
    .S0(net406),
    .S1(net395),
    .X(_2271_));
 sky130_fd_sc_hd__mux4_1 _4715_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ),
    .S0(net405),
    .S1(net395),
    .X(_2272_));
 sky130_fd_sc_hd__mux2_1 _4716_ (.A0(_2272_),
    .A1(_2271_),
    .S(net386),
    .X(_2273_));
 sky130_fd_sc_hd__mux2_1 _4717_ (.A0(_2273_),
    .A1(_2270_),
    .S(net382),
    .X(_0000_));
 sky130_fd_sc_hd__mux4_1 _4718_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ),
    .S0(net405),
    .S1(net395),
    .X(_2274_));
 sky130_fd_sc_hd__mux4_1 _4719_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ),
    .S0(net405),
    .S1(net395),
    .X(_2275_));
 sky130_fd_sc_hd__mux2_1 _4720_ (.A0(_2274_),
    .A1(_2275_),
    .S(net386),
    .X(_2276_));
 sky130_fd_sc_hd__mux4_1 _4721_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ),
    .S0(net405),
    .S1(net395),
    .X(_2277_));
 sky130_fd_sc_hd__mux4_1 _4722_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ),
    .S0(net405),
    .S1(net395),
    .X(_2278_));
 sky130_fd_sc_hd__mux2_1 _4723_ (.A0(_2278_),
    .A1(_2277_),
    .S(net386),
    .X(_2279_));
 sky130_fd_sc_hd__mux2_1 _4724_ (.A0(_2279_),
    .A1(_2276_),
    .S(net383),
    .X(_0011_));
 sky130_fd_sc_hd__mux4_1 _4725_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ),
    .S0(net405),
    .S1(net395),
    .X(_2280_));
 sky130_fd_sc_hd__mux4_1 _4726_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ),
    .S0(net405),
    .S1(net395),
    .X(_2281_));
 sky130_fd_sc_hd__mux2_1 _4727_ (.A0(_2280_),
    .A1(_2281_),
    .S(net386),
    .X(_2282_));
 sky130_fd_sc_hd__mux4_1 _4728_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ),
    .S0(net405),
    .S1(net395),
    .X(_2283_));
 sky130_fd_sc_hd__mux4_1 _4729_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ),
    .S0(net406),
    .S1(net395),
    .X(_2284_));
 sky130_fd_sc_hd__mux2_1 _4730_ (.A0(_2284_),
    .A1(_2283_),
    .S(net386),
    .X(_2285_));
 sky130_fd_sc_hd__mux2_1 _4731_ (.A0(_2285_),
    .A1(_2282_),
    .S(net382),
    .X(_0022_));
 sky130_fd_sc_hd__mux4_1 _4732_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ),
    .S0(net405),
    .S1(net395),
    .X(_2286_));
 sky130_fd_sc_hd__mux4_1 _4733_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ),
    .S0(net405),
    .S1(net395),
    .X(_2287_));
 sky130_fd_sc_hd__mux2_1 _4734_ (.A0(_2286_),
    .A1(_2287_),
    .S(net386),
    .X(_2288_));
 sky130_fd_sc_hd__mux4_1 _4735_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ),
    .S0(net405),
    .S1(net395),
    .X(_2289_));
 sky130_fd_sc_hd__mux4_1 _4736_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ),
    .S0(net405),
    .S1(net395),
    .X(_2290_));
 sky130_fd_sc_hd__mux2_1 _4737_ (.A0(_2290_),
    .A1(_2289_),
    .S(net387),
    .X(_2291_));
 sky130_fd_sc_hd__mux2_1 _4738_ (.A0(_2291_),
    .A1(_2288_),
    .S(net383),
    .X(_0025_));
 sky130_fd_sc_hd__mux4_1 _4739_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ),
    .S0(net408),
    .S1(net398),
    .X(_2292_));
 sky130_fd_sc_hd__mux4_1 _4740_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ),
    .S0(net408),
    .S1(net398),
    .X(_2293_));
 sky130_fd_sc_hd__mux2_1 _4741_ (.A0(_2292_),
    .A1(_2293_),
    .S(net388),
    .X(_2294_));
 sky130_fd_sc_hd__mux4_1 _4742_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ),
    .S0(net406),
    .S1(net396),
    .X(_2295_));
 sky130_fd_sc_hd__mux4_1 _4743_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ),
    .S0(net406),
    .S1(net396),
    .X(_2296_));
 sky130_fd_sc_hd__mux2_1 _4744_ (.A0(_2296_),
    .A1(_2295_),
    .S(net386),
    .X(_2297_));
 sky130_fd_sc_hd__mux2_1 _4745_ (.A0(_2297_),
    .A1(_2294_),
    .S(net382),
    .X(_0026_));
 sky130_fd_sc_hd__mux4_1 _4746_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ),
    .S0(net404),
    .S1(net394),
    .X(_2298_));
 sky130_fd_sc_hd__mux4_1 _4747_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ),
    .S0(net404),
    .S1(net397),
    .X(_2299_));
 sky130_fd_sc_hd__mux2_1 _4748_ (.A0(_2298_),
    .A1(_2299_),
    .S(net387),
    .X(_2300_));
 sky130_fd_sc_hd__mux4_1 _4749_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ),
    .S0(net404),
    .S1(net394),
    .X(_2301_));
 sky130_fd_sc_hd__mux4_1 _4750_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ),
    .S0(net407),
    .S1(net394),
    .X(_2302_));
 sky130_fd_sc_hd__mux2_1 _4751_ (.A0(_2302_),
    .A1(_2301_),
    .S(net387),
    .X(_2303_));
 sky130_fd_sc_hd__mux2_1 _4752_ (.A0(_2303_),
    .A1(_2300_),
    .S(net382),
    .X(_0027_));
 sky130_fd_sc_hd__mux4_1 _4753_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ),
    .S0(net403),
    .S1(net393),
    .X(_2304_));
 sky130_fd_sc_hd__mux4_1 _4754_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ),
    .S0(net403),
    .S1(net393),
    .X(_2305_));
 sky130_fd_sc_hd__mux2_1 _4755_ (.A0(_2304_),
    .A1(_2305_),
    .S(net388),
    .X(_2306_));
 sky130_fd_sc_hd__mux4_1 _4756_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ),
    .S0(net403),
    .S1(net393),
    .X(_2307_));
 sky130_fd_sc_hd__mux4_1 _4757_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ),
    .S0(net403),
    .S1(net393),
    .X(_2308_));
 sky130_fd_sc_hd__mux2_1 _4758_ (.A0(_2308_),
    .A1(_2307_),
    .S(net388),
    .X(_2309_));
 sky130_fd_sc_hd__mux2_1 _4759_ (.A0(_2309_),
    .A1(_2306_),
    .S(net382),
    .X(_0028_));
 sky130_fd_sc_hd__mux4_1 _4760_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ),
    .S0(net399),
    .S1(net389),
    .X(_2310_));
 sky130_fd_sc_hd__mux4_1 _4761_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ),
    .S0(net400),
    .S1(net390),
    .X(_2311_));
 sky130_fd_sc_hd__mux2_1 _4762_ (.A0(_2310_),
    .A1(_2311_),
    .S(net384),
    .X(_2312_));
 sky130_fd_sc_hd__mux4_1 _4763_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ),
    .S0(net400),
    .S1(net390),
    .X(_2313_));
 sky130_fd_sc_hd__mux4_1 _4764_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ),
    .S0(net400),
    .S1(net390),
    .X(_2314_));
 sky130_fd_sc_hd__mux2_1 _4765_ (.A0(_2314_),
    .A1(_2313_),
    .S(net384),
    .X(_2315_));
 sky130_fd_sc_hd__mux2_1 _4766_ (.A0(_2315_),
    .A1(_2312_),
    .S(net381),
    .X(_0029_));
 sky130_fd_sc_hd__mux4_1 _4767_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ),
    .S0(net400),
    .S1(net390),
    .X(_2316_));
 sky130_fd_sc_hd__mux4_1 _4768_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ),
    .S0(net400),
    .S1(net390),
    .X(_2317_));
 sky130_fd_sc_hd__mux2_1 _4769_ (.A0(_2316_),
    .A1(_2317_),
    .S(net384),
    .X(_2318_));
 sky130_fd_sc_hd__mux4_1 _4770_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ),
    .S1(net398),
    .X(_2319_));
 sky130_fd_sc_hd__mux4_1 _4771_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ),
    .S0(net402),
    .S1(net392),
    .X(_2320_));
 sky130_fd_sc_hd__mux2_1 _4772_ (.A0(_2320_),
    .A1(_2319_),
    .S(net385),
    .X(_2321_));
 sky130_fd_sc_hd__mux2_1 _4773_ (.A0(_2321_),
    .A1(_2318_),
    .S(net381),
    .X(_0030_));
 sky130_fd_sc_hd__mux4_1 _4774_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ),
    .S0(net403),
    .S1(net393),
    .X(_2322_));
 sky130_fd_sc_hd__mux4_1 _4775_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ),
    .S0(net408),
    .S1(net393),
    .X(_2323_));
 sky130_fd_sc_hd__mux2_1 _4776_ (.A0(_2322_),
    .A1(_2323_),
    .S(net388),
    .X(_2324_));
 sky130_fd_sc_hd__mux4_1 _4777_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ),
    .S0(net403),
    .S1(net393),
    .X(_2325_));
 sky130_fd_sc_hd__mux4_1 _4778_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ),
    .S0(net403),
    .S1(net393),
    .X(_2326_));
 sky130_fd_sc_hd__mux2_1 _4779_ (.A0(_2326_),
    .A1(_2325_),
    .S(net388),
    .X(_2327_));
 sky130_fd_sc_hd__mux2_1 _4780_ (.A0(_2327_),
    .A1(_2324_),
    .S(net382),
    .X(_0031_));
 sky130_fd_sc_hd__mux4_1 _4781_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ),
    .S1(net398),
    .X(_2328_));
 sky130_fd_sc_hd__mux4_1 _4782_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ),
    .S1(net398),
    .X(_2329_));
 sky130_fd_sc_hd__mux2_1 _4783_ (.A0(_2328_),
    .A1(_2329_),
    .S(net385),
    .X(_2330_));
 sky130_fd_sc_hd__mux4_1 _4784_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ),
    .S0(net402),
    .S1(net392),
    .X(_2331_));
 sky130_fd_sc_hd__mux4_1 _4785_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ),
    .S0(net402),
    .S1(net398),
    .X(_2332_));
 sky130_fd_sc_hd__mux2_1 _4786_ (.A0(_2332_),
    .A1(_2331_),
    .S(net385),
    .X(_2333_));
 sky130_fd_sc_hd__mux2_1 _4787_ (.A0(_2333_),
    .A1(_2330_),
    .S(net383),
    .X(_0001_));
 sky130_fd_sc_hd__mux4_1 _4788_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ),
    .S0(net400),
    .S1(net390),
    .X(_2334_));
 sky130_fd_sc_hd__mux4_1 _4789_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ),
    .S0(net400),
    .S1(net390),
    .X(_2335_));
 sky130_fd_sc_hd__mux2_1 _4790_ (.A0(_2334_),
    .A1(_2335_),
    .S(net384),
    .X(_2336_));
 sky130_fd_sc_hd__mux4_1 _4791_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ),
    .S0(net400),
    .S1(net390),
    .X(_2337_));
 sky130_fd_sc_hd__mux4_1 _4792_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ),
    .S0(net400),
    .S1(net390),
    .X(_2338_));
 sky130_fd_sc_hd__mux2_1 _4793_ (.A0(_2338_),
    .A1(_2337_),
    .S(net384),
    .X(_2339_));
 sky130_fd_sc_hd__mux2_1 _4794_ (.A0(_2339_),
    .A1(_2336_),
    .S(net381),
    .X(_0002_));
 sky130_fd_sc_hd__mux4_1 _4795_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ),
    .S0(net403),
    .S1(net393),
    .X(_2340_));
 sky130_fd_sc_hd__mux4_1 _4796_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ),
    .S0(net406),
    .S1(net396),
    .X(_2341_));
 sky130_fd_sc_hd__mux2_1 _4797_ (.A0(_2340_),
    .A1(_2341_),
    .S(net386),
    .X(_2342_));
 sky130_fd_sc_hd__mux4_1 _4798_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ),
    .S0(net403),
    .S1(net398),
    .X(_2343_));
 sky130_fd_sc_hd__mux4_1 _4799_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ),
    .S0(net403),
    .S1(net398),
    .X(_2344_));
 sky130_fd_sc_hd__mux2_1 _4800_ (.A0(_2344_),
    .A1(_2343_),
    .S(net388),
    .X(_2345_));
 sky130_fd_sc_hd__mux2_1 _4801_ (.A0(_2345_),
    .A1(_2342_),
    .S(net382),
    .X(_0003_));
 sky130_fd_sc_hd__mux4_1 _4802_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ),
    .S0(net403),
    .S1(net393),
    .X(_2346_));
 sky130_fd_sc_hd__mux4_1 _4803_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ),
    .S0(net406),
    .S1(net396),
    .X(_2347_));
 sky130_fd_sc_hd__mux2_1 _4804_ (.A0(_2346_),
    .A1(_2347_),
    .S(net386),
    .X(_2348_));
 sky130_fd_sc_hd__mux4_1 _4805_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ),
    .S0(net406),
    .S1(net396),
    .X(_2349_));
 sky130_fd_sc_hd__mux4_1 _4806_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ),
    .S0(net403),
    .S1(net393),
    .X(_2350_));
 sky130_fd_sc_hd__mux2_1 _4807_ (.A0(_2350_),
    .A1(_2349_),
    .S(net386),
    .X(_2351_));
 sky130_fd_sc_hd__mux2_1 _4808_ (.A0(_2351_),
    .A1(_2348_),
    .S(net383),
    .X(_0004_));
 sky130_fd_sc_hd__mux4_1 _4809_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ),
    .S0(net407),
    .S1(net397),
    .X(_2352_));
 sky130_fd_sc_hd__mux4_1 _4810_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ),
    .S0(net404),
    .S1(net397),
    .X(_2353_));
 sky130_fd_sc_hd__mux2_1 _4811_ (.A0(_2352_),
    .A1(_2353_),
    .S(net387),
    .X(_2354_));
 sky130_fd_sc_hd__mux4_1 _4812_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ),
    .S0(net407),
    .S1(net397),
    .X(_2355_));
 sky130_fd_sc_hd__mux4_1 _4813_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ),
    .S0(net407),
    .S1(net397),
    .X(_2356_));
 sky130_fd_sc_hd__mux2_1 _4814_ (.A0(_2356_),
    .A1(_2355_),
    .S(net387),
    .X(_2357_));
 sky130_fd_sc_hd__mux2_1 _4815_ (.A0(_2357_),
    .A1(_2354_),
    .S(net383),
    .X(_0005_));
 sky130_fd_sc_hd__mux4_1 _4816_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ),
    .S0(net404),
    .S1(net394),
    .X(_2358_));
 sky130_fd_sc_hd__mux4_1 _4817_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ),
    .S0(net404),
    .S1(net394),
    .X(_2359_));
 sky130_fd_sc_hd__mux2_1 _4818_ (.A0(_2358_),
    .A1(_2359_),
    .S(net387),
    .X(_2360_));
 sky130_fd_sc_hd__mux4_1 _4819_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ),
    .S0(net404),
    .S1(net394),
    .X(_2361_));
 sky130_fd_sc_hd__mux4_1 _4820_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ),
    .S0(net404),
    .S1(net394),
    .X(_2362_));
 sky130_fd_sc_hd__mux2_1 _4821_ (.A0(_2362_),
    .A1(_2361_),
    .S(net387),
    .X(_2363_));
 sky130_fd_sc_hd__mux2_1 _4822_ (.A0(_2363_),
    .A1(_2360_),
    .S(net382),
    .X(_0006_));
 sky130_fd_sc_hd__mux4_1 _4823_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ),
    .S0(net402),
    .S1(net392),
    .X(_2364_));
 sky130_fd_sc_hd__mux4_1 _4824_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ),
    .S0(net402),
    .S1(net392),
    .X(_2365_));
 sky130_fd_sc_hd__mux2_1 _4825_ (.A0(_2364_),
    .A1(_2365_),
    .S(net385),
    .X(_2366_));
 sky130_fd_sc_hd__mux4_1 _4826_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ),
    .S0(net402),
    .S1(net392),
    .X(_2367_));
 sky130_fd_sc_hd__mux4_1 _4827_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ),
    .S0(net402),
    .S1(net392),
    .X(_2368_));
 sky130_fd_sc_hd__mux2_1 _4828_ (.A0(_2368_),
    .A1(_2367_),
    .S(net385),
    .X(_2369_));
 sky130_fd_sc_hd__mux2_1 _4829_ (.A0(_2369_),
    .A1(_2366_),
    .S(net381),
    .X(_0007_));
 sky130_fd_sc_hd__mux4_1 _4830_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ),
    .S0(net403),
    .S1(net393),
    .X(_2370_));
 sky130_fd_sc_hd__mux4_1 _4831_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ),
    .S0(net408),
    .S1(net393),
    .X(_2371_));
 sky130_fd_sc_hd__mux2_1 _4832_ (.A0(_2370_),
    .A1(_2371_),
    .S(net388),
    .X(_2372_));
 sky130_fd_sc_hd__mux4_1 _4833_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ),
    .S0(net403),
    .S1(net393),
    .X(_2373_));
 sky130_fd_sc_hd__mux4_1 _4834_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ),
    .S0(net402),
    .S1(net392),
    .X(_2374_));
 sky130_fd_sc_hd__mux2_1 _4835_ (.A0(_2374_),
    .A1(_2373_),
    .S(net388),
    .X(_2375_));
 sky130_fd_sc_hd__mux2_1 _4836_ (.A0(_2375_),
    .A1(_2372_),
    .S(net382),
    .X(_0008_));
 sky130_fd_sc_hd__mux4_1 _4837_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ),
    .S0(net407),
    .S1(net394),
    .X(_2376_));
 sky130_fd_sc_hd__mux4_1 _4838_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ),
    .S0(net407),
    .S1(net397),
    .X(_2377_));
 sky130_fd_sc_hd__mux2_1 _4839_ (.A0(_2376_),
    .A1(_2377_),
    .S(net387),
    .X(_2378_));
 sky130_fd_sc_hd__mux4_1 _4840_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ),
    .S0(net407),
    .S1(net394),
    .X(_2379_));
 sky130_fd_sc_hd__mux4_1 _4841_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ),
    .S0(net404),
    .S1(net394),
    .X(_2380_));
 sky130_fd_sc_hd__mux2_1 _4842_ (.A0(_2380_),
    .A1(_2379_),
    .S(net387),
    .X(_2381_));
 sky130_fd_sc_hd__mux2_1 _4843_ (.A0(_2381_),
    .A1(_2378_),
    .S(net382),
    .X(_0009_));
 sky130_fd_sc_hd__mux4_1 _4844_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ),
    .S0(net404),
    .S1(net394),
    .X(_2382_));
 sky130_fd_sc_hd__mux4_1 _4845_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ),
    .S0(net404),
    .S1(net394),
    .X(_2383_));
 sky130_fd_sc_hd__mux2_1 _4846_ (.A0(_2382_),
    .A1(_2383_),
    .S(net387),
    .X(_2384_));
 sky130_fd_sc_hd__mux4_1 _4847_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ),
    .S0(net404),
    .S1(net394),
    .X(_2385_));
 sky130_fd_sc_hd__mux4_1 _4848_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ),
    .S0(net404),
    .S1(net394),
    .X(_2386_));
 sky130_fd_sc_hd__mux2_1 _4849_ (.A0(_2386_),
    .A1(_2385_),
    .S(net387),
    .X(_2387_));
 sky130_fd_sc_hd__mux2_1 _4850_ (.A0(_2387_),
    .A1(_2384_),
    .S(net382),
    .X(_0010_));
 sky130_fd_sc_hd__mux4_1 _4851_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ),
    .S0(net401),
    .S1(net391),
    .X(_2388_));
 sky130_fd_sc_hd__mux4_1 _4852_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ),
    .S0(net401),
    .S1(net391),
    .X(_2389_));
 sky130_fd_sc_hd__mux2_1 _4853_ (.A0(_2388_),
    .A1(_2389_),
    .S(net385),
    .X(_2390_));
 sky130_fd_sc_hd__mux4_1 _4854_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ),
    .S0(net401),
    .S1(net391),
    .X(_2391_));
 sky130_fd_sc_hd__mux4_1 _4855_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ),
    .S0(net401),
    .S1(net391),
    .X(_2392_));
 sky130_fd_sc_hd__mux2_1 _4856_ (.A0(_2392_),
    .A1(_2391_),
    .S(net385),
    .X(_2393_));
 sky130_fd_sc_hd__mux2_1 _4857_ (.A0(_2393_),
    .A1(_2390_),
    .S(net381),
    .X(_0012_));
 sky130_fd_sc_hd__mux4_1 _4858_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ),
    .S0(net401),
    .S1(net391),
    .X(_2394_));
 sky130_fd_sc_hd__mux4_1 _4859_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ),
    .S0(net401),
    .S1(net391),
    .X(_2395_));
 sky130_fd_sc_hd__mux2_1 _4860_ (.A0(_2394_),
    .A1(_2395_),
    .S(net384),
    .X(_2396_));
 sky130_fd_sc_hd__mux4_1 _4861_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ),
    .S0(net401),
    .S1(net391),
    .X(_2397_));
 sky130_fd_sc_hd__mux4_1 _4862_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ),
    .S0(net401),
    .S1(net391),
    .X(_2398_));
 sky130_fd_sc_hd__mux2_1 _4863_ (.A0(_2398_),
    .A1(_2397_),
    .S(net384),
    .X(_2399_));
 sky130_fd_sc_hd__mux2_1 _4864_ (.A0(_2399_),
    .A1(_2396_),
    .S(net381),
    .X(_0013_));
 sky130_fd_sc_hd__mux4_1 _4865_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ),
    .S0(net405),
    .S1(net396),
    .X(_2400_));
 sky130_fd_sc_hd__mux4_1 _4866_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ),
    .S0(net406),
    .S1(net396),
    .X(_2401_));
 sky130_fd_sc_hd__mux2_1 _4867_ (.A0(_2400_),
    .A1(_2401_),
    .S(net386),
    .X(_2402_));
 sky130_fd_sc_hd__mux4_1 _4868_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ),
    .S0(net406),
    .S1(net396),
    .X(_2403_));
 sky130_fd_sc_hd__mux4_1 _4869_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ),
    .S0(net406),
    .S1(net396),
    .X(_2404_));
 sky130_fd_sc_hd__mux2_1 _4870_ (.A0(_2404_),
    .A1(_2403_),
    .S(net386),
    .X(_2405_));
 sky130_fd_sc_hd__mux2_1 _4871_ (.A0(_2405_),
    .A1(_2402_),
    .S(net383),
    .X(_0014_));
 sky130_fd_sc_hd__mux4_1 _4872_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ),
    .S0(net401),
    .S1(net391),
    .X(_2406_));
 sky130_fd_sc_hd__mux4_1 _4873_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ),
    .S0(net400),
    .S1(net390),
    .X(_2407_));
 sky130_fd_sc_hd__mux2_1 _4874_ (.A0(_2406_),
    .A1(_2407_),
    .S(net385),
    .X(_2408_));
 sky130_fd_sc_hd__mux4_1 _4875_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ),
    .S0(net401),
    .S1(net391),
    .X(_2409_));
 sky130_fd_sc_hd__mux4_1 _4876_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ),
    .S0(net401),
    .S1(net391),
    .X(_2410_));
 sky130_fd_sc_hd__mux2_1 _4877_ (.A0(_2410_),
    .A1(_2409_),
    .S(net385),
    .X(_2411_));
 sky130_fd_sc_hd__mux2_1 _4878_ (.A0(_2411_),
    .A1(_2408_),
    .S(net381),
    .X(_0015_));
 sky130_fd_sc_hd__mux4_1 _4879_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ),
    .S0(net406),
    .S1(net396),
    .X(_2412_));
 sky130_fd_sc_hd__mux4_1 _4880_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ),
    .S0(net406),
    .S1(net396),
    .X(_2413_));
 sky130_fd_sc_hd__mux2_1 _4881_ (.A0(_2412_),
    .A1(_2413_),
    .S(net386),
    .X(_2414_));
 sky130_fd_sc_hd__mux4_1 _4882_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ),
    .S0(net406),
    .S1(net396),
    .X(_2415_));
 sky130_fd_sc_hd__mux4_1 _4883_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ),
    .S0(net406),
    .S1(net396),
    .X(_2416_));
 sky130_fd_sc_hd__mux2_1 _4884_ (.A0(_2416_),
    .A1(_2415_),
    .S(net386),
    .X(_2417_));
 sky130_fd_sc_hd__mux2_1 _4885_ (.A0(_2417_),
    .A1(_2414_),
    .S(net382),
    .X(_0016_));
 sky130_fd_sc_hd__mux4_1 _4886_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ),
    .S0(net399),
    .S1(net389),
    .X(_2418_));
 sky130_fd_sc_hd__mux4_1 _4887_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ),
    .S0(net399),
    .S1(net389),
    .X(_2419_));
 sky130_fd_sc_hd__mux2_1 _4888_ (.A0(_2418_),
    .A1(_2419_),
    .S(net384),
    .X(_2420_));
 sky130_fd_sc_hd__mux4_1 _4889_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ),
    .S0(net399),
    .S1(net389),
    .X(_2421_));
 sky130_fd_sc_hd__mux4_1 _4890_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ),
    .S0(net399),
    .S1(net389),
    .X(_2422_));
 sky130_fd_sc_hd__mux2_1 _4891_ (.A0(_2422_),
    .A1(_2421_),
    .S(net384),
    .X(_2423_));
 sky130_fd_sc_hd__mux2_1 _4892_ (.A0(_2423_),
    .A1(_2420_),
    .S(net381),
    .X(_0017_));
 sky130_fd_sc_hd__mux4_1 _4893_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ),
    .S0(net401),
    .S1(net391),
    .X(_2424_));
 sky130_fd_sc_hd__mux4_1 _4894_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ),
    .S0(net401),
    .S1(net391),
    .X(_2425_));
 sky130_fd_sc_hd__mux2_1 _4895_ (.A0(_2424_),
    .A1(_2425_),
    .S(net384),
    .X(_2426_));
 sky130_fd_sc_hd__mux4_1 _4896_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ),
    .S0(net401),
    .S1(net391),
    .X(_2427_));
 sky130_fd_sc_hd__mux4_1 _4897_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ),
    .S0(net401),
    .S1(net391),
    .X(_2428_));
 sky130_fd_sc_hd__mux2_1 _4898_ (.A0(_2428_),
    .A1(_2427_),
    .S(net385),
    .X(_2429_));
 sky130_fd_sc_hd__mux2_1 _4899_ (.A0(_2429_),
    .A1(_2426_),
    .S(net381),
    .X(_0018_));
 sky130_fd_sc_hd__mux4_1 _4900_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ),
    .S0(net403),
    .S1(net393),
    .X(_2430_));
 sky130_fd_sc_hd__mux4_1 _4901_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ),
    .S0(net402),
    .S1(net392),
    .X(_2431_));
 sky130_fd_sc_hd__mux2_1 _4902_ (.A0(_2430_),
    .A1(_2431_),
    .S(net385),
    .X(_2432_));
 sky130_fd_sc_hd__mux4_1 _4903_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ),
    .S0(net402),
    .S1(net392),
    .X(_2433_));
 sky130_fd_sc_hd__mux4_1 _4904_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ),
    .S0(net403),
    .S1(net393),
    .X(_2434_));
 sky130_fd_sc_hd__mux2_1 _4905_ (.A0(_2434_),
    .A1(_2433_),
    .S(net385),
    .X(_2435_));
 sky130_fd_sc_hd__mux2_1 _4906_ (.A0(_2435_),
    .A1(_2432_),
    .S(net381),
    .X(_0019_));
 sky130_fd_sc_hd__mux4_1 _4907_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ),
    .S0(net399),
    .S1(net389),
    .X(_2436_));
 sky130_fd_sc_hd__mux4_1 _4908_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ),
    .S0(net399),
    .S1(net389),
    .X(_2437_));
 sky130_fd_sc_hd__mux2_1 _4909_ (.A0(_2436_),
    .A1(_2437_),
    .S(net384),
    .X(_2438_));
 sky130_fd_sc_hd__mux4_1 _4910_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ),
    .S0(net399),
    .S1(net389),
    .X(_2439_));
 sky130_fd_sc_hd__mux4_1 _4911_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ),
    .S0(net399),
    .S1(net389),
    .X(_2440_));
 sky130_fd_sc_hd__mux2_1 _4912_ (.A0(_2440_),
    .A1(_2439_),
    .S(net384),
    .X(_2441_));
 sky130_fd_sc_hd__mux2_1 _4913_ (.A0(_2441_),
    .A1(_2438_),
    .S(net381),
    .X(_0020_));
 sky130_fd_sc_hd__mux4_1 _4914_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ),
    .S0(net399),
    .S1(net390),
    .X(_2442_));
 sky130_fd_sc_hd__mux4_1 _4915_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ),
    .S0(net400),
    .S1(net389),
    .X(_2443_));
 sky130_fd_sc_hd__mux2_1 _4916_ (.A0(_2442_),
    .A1(_2443_),
    .S(net384),
    .X(_2444_));
 sky130_fd_sc_hd__mux4_1 _4917_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ),
    .S0(net399),
    .S1(net389),
    .X(_2445_));
 sky130_fd_sc_hd__mux4_1 _4918_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ),
    .S0(net399),
    .S1(net389),
    .X(_2446_));
 sky130_fd_sc_hd__mux2_1 _4919_ (.A0(_2446_),
    .A1(_2445_),
    .S(net384),
    .X(_2447_));
 sky130_fd_sc_hd__mux2_1 _4920_ (.A0(_2447_),
    .A1(_2444_),
    .S(net381),
    .X(_0021_));
 sky130_fd_sc_hd__mux4_1 _4921_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ),
    .S0(net399),
    .S1(net389),
    .X(_2448_));
 sky130_fd_sc_hd__mux4_1 _4922_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ),
    .S0(net399),
    .S1(net389),
    .X(_2449_));
 sky130_fd_sc_hd__mux2_1 _4923_ (.A0(_2448_),
    .A1(_2449_),
    .S(net384),
    .X(_2450_));
 sky130_fd_sc_hd__mux4_1 _4924_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ),
    .S0(net399),
    .S1(net389),
    .X(_2451_));
 sky130_fd_sc_hd__mux4_1 _4925_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ),
    .S0(net399),
    .S1(net389),
    .X(_2452_));
 sky130_fd_sc_hd__mux2_1 _4926_ (.A0(_2452_),
    .A1(_2451_),
    .S(net384),
    .X(_2453_));
 sky130_fd_sc_hd__mux2_1 _4927_ (.A0(_2453_),
    .A1(_2450_),
    .S(net381),
    .X(_0023_));
 sky130_fd_sc_hd__mux4_1 _4928_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ),
    .S0(net402),
    .S1(net392),
    .X(_2454_));
 sky130_fd_sc_hd__mux4_1 _4929_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ),
    .S0(net402),
    .S1(net392),
    .X(_2455_));
 sky130_fd_sc_hd__mux2_1 _4930_ (.A0(_2454_),
    .A1(_2455_),
    .S(net385),
    .X(_2456_));
 sky130_fd_sc_hd__mux4_1 _4931_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ),
    .S0(net401),
    .S1(net392),
    .X(_2457_));
 sky130_fd_sc_hd__mux4_1 _4932_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ),
    .S0(net402),
    .S1(net391),
    .X(_2458_));
 sky130_fd_sc_hd__mux2_1 _4933_ (.A0(_2458_),
    .A1(_2457_),
    .S(net385),
    .X(_2459_));
 sky130_fd_sc_hd__mux2_1 _4934_ (.A0(_2459_),
    .A1(_2456_),
    .S(net381),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _4935_ (.A(net462),
    .B(net2133),
    .X(_0069_));
 sky130_fd_sc_hd__nor2_1 _4936_ (.A(net479),
    .B(net1508),
    .Y(_0080_));
 sky130_fd_sc_hd__and2_1 _4937_ (.A(net467),
    .B(net1780),
    .X(_0091_));
 sky130_fd_sc_hd__and2_1 _4938_ (.A(net464),
    .B(net2135),
    .X(_0094_));
 sky130_fd_sc_hd__and2_1 _4939_ (.A(net458),
    .B(net2127),
    .X(_0095_));
 sky130_fd_sc_hd__and2_1 _4940_ (.A(net458),
    .B(net2035),
    .X(_0096_));
 sky130_fd_sc_hd__and2_1 _4941_ (.A(net453),
    .B(net2159),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _4942_ (.A(net446),
    .B(net2054),
    .X(_0098_));
 sky130_fd_sc_hd__and2_1 _4943_ (.A(net447),
    .B(net2139),
    .X(_0099_));
 sky130_fd_sc_hd__and2_1 _4944_ (.A(net461),
    .B(net1919),
    .X(_0100_));
 sky130_fd_sc_hd__and2_1 _4945_ (.A(net449),
    .B(net2066),
    .X(_0070_));
 sky130_fd_sc_hd__and2_1 _4946_ (.A(net447),
    .B(net2009),
    .X(_0071_));
 sky130_fd_sc_hd__and2_1 _4947_ (.A(net461),
    .B(net1822),
    .X(_0072_));
 sky130_fd_sc_hd__and2_1 _4948_ (.A(net462),
    .B(net2091),
    .X(_0073_));
 sky130_fd_sc_hd__and2_1 _4949_ (.A(net458),
    .B(net2025),
    .X(_0074_));
 sky130_fd_sc_hd__and2_1 _4950_ (.A(net457),
    .B(net1709),
    .X(_0075_));
 sky130_fd_sc_hd__and2_1 _4951_ (.A(net453),
    .B(net2122),
    .X(_0076_));
 sky130_fd_sc_hd__and2_1 _4952_ (.A(net453),
    .B(net2067),
    .X(_0077_));
 sky130_fd_sc_hd__and2_1 _4953_ (.A(net471),
    .B(net1892),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _4954_ (.A(net458),
    .B(net767),
    .X(_0079_));
 sky130_fd_sc_hd__and2_1 _4955_ (.A(net446),
    .B(net2140),
    .X(_0081_));
 sky130_fd_sc_hd__and2_1 _4956_ (.A(net445),
    .B(net1963),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _4957_ (.A(net467),
    .B(net1988),
    .X(_0083_));
 sky130_fd_sc_hd__and2_1 _4958_ (.A(net446),
    .B(net2065),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _4959_ (.A(net461),
    .B(net863),
    .X(_0085_));
 sky130_fd_sc_hd__and2_1 _4960_ (.A(net446),
    .B(net2153),
    .X(_0086_));
 sky130_fd_sc_hd__and2_1 _4961_ (.A(net445),
    .B(net1993),
    .X(_0087_));
 sky130_fd_sc_hd__and2_1 _4962_ (.A(net451),
    .B(net1991),
    .X(_0088_));
 sky130_fd_sc_hd__and2_1 _4963_ (.A(net441),
    .B(net1968),
    .X(_0089_));
 sky130_fd_sc_hd__and2_1 _4964_ (.A(net442),
    .B(net2062),
    .X(_0090_));
 sky130_fd_sc_hd__and2_1 _4965_ (.A(net447),
    .B(net1992),
    .X(_0092_));
 sky130_fd_sc_hd__and2_1 _4966_ (.A(net451),
    .B(net623),
    .X(_0093_));
 sky130_fd_sc_hd__mux4_1 _4967_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ),
    .S0(net434),
    .S1(net423),
    .X(_2460_));
 sky130_fd_sc_hd__mux4_1 _4968_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ),
    .S0(net434),
    .S1(net423),
    .X(_2461_));
 sky130_fd_sc_hd__mux2_1 _4969_ (.A0(_2460_),
    .A1(_2461_),
    .S(net415),
    .X(_2462_));
 sky130_fd_sc_hd__mux4_1 _4970_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ),
    .S0(net435),
    .S1(net423),
    .X(_2463_));
 sky130_fd_sc_hd__mux4_1 _4971_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ),
    .S0(net434),
    .S1(net423),
    .X(_2464_));
 sky130_fd_sc_hd__mux2_1 _4972_ (.A0(_2464_),
    .A1(_2463_),
    .S(net415),
    .X(_2465_));
 sky130_fd_sc_hd__mux2_1 _4973_ (.A0(_2465_),
    .A1(_2462_),
    .S(net409),
    .X(_0032_));
 sky130_fd_sc_hd__mux4_1 _4974_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ),
    .S0(net435),
    .S1(net423),
    .X(_2466_));
 sky130_fd_sc_hd__mux4_1 _4975_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ),
    .S0(net435),
    .S1(net423),
    .X(_2467_));
 sky130_fd_sc_hd__mux2_1 _4976_ (.A0(_2466_),
    .A1(_2467_),
    .S(net415),
    .X(_2468_));
 sky130_fd_sc_hd__mux4_1 _4977_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ),
    .S0(net435),
    .S1(net423),
    .X(_2469_));
 sky130_fd_sc_hd__mux4_1 _4978_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ),
    .S0(net435),
    .S1(net423),
    .X(_2470_));
 sky130_fd_sc_hd__mux2_1 _4979_ (.A0(_2470_),
    .A1(_2469_),
    .S(net415),
    .X(_2471_));
 sky130_fd_sc_hd__mux2_1 _4980_ (.A0(_2471_),
    .A1(_2468_),
    .S(net409),
    .X(_0043_));
 sky130_fd_sc_hd__mux4_1 _4981_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ),
    .S0(net435),
    .S1(net423),
    .X(_2472_));
 sky130_fd_sc_hd__mux4_1 _4982_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ),
    .S0(net435),
    .S1(net423),
    .X(_2473_));
 sky130_fd_sc_hd__mux2_1 _4983_ (.A0(_2472_),
    .A1(_2473_),
    .S(net415),
    .X(_2474_));
 sky130_fd_sc_hd__mux4_1 _4984_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ),
    .S0(net435),
    .S1(net423),
    .X(_2475_));
 sky130_fd_sc_hd__mux4_1 _4985_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ),
    .S0(net435),
    .S1(net423),
    .X(_2476_));
 sky130_fd_sc_hd__mux2_1 _4986_ (.A0(_2476_),
    .A1(_2475_),
    .S(net415),
    .X(_2477_));
 sky130_fd_sc_hd__mux2_1 _4987_ (.A0(_2477_),
    .A1(_2474_),
    .S(net409),
    .X(_0054_));
 sky130_fd_sc_hd__mux4_1 _4988_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ),
    .S0(net434),
    .S1(net423),
    .X(_2478_));
 sky130_fd_sc_hd__mux4_1 _4989_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ),
    .S0(net435),
    .S1(net423),
    .X(_2479_));
 sky130_fd_sc_hd__mux2_1 _4990_ (.A0(_2478_),
    .A1(_2479_),
    .S(net415),
    .X(_2480_));
 sky130_fd_sc_hd__mux4_1 _4991_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ),
    .S0(net434),
    .S1(net423),
    .X(_2481_));
 sky130_fd_sc_hd__mux4_1 _4992_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ),
    .S0(net435),
    .S1(net423),
    .X(_2482_));
 sky130_fd_sc_hd__mux2_1 _4993_ (.A0(_2482_),
    .A1(_2481_),
    .S(net415),
    .X(_2483_));
 sky130_fd_sc_hd__mux2_1 _4994_ (.A0(_2483_),
    .A1(_2480_),
    .S(net409),
    .X(_0057_));
 sky130_fd_sc_hd__mux4_1 _4995_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ),
    .S0(net432),
    .S1(net426),
    .X(_2484_));
 sky130_fd_sc_hd__mux4_1 _4996_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ),
    .S0(net432),
    .S1(net426),
    .X(_2485_));
 sky130_fd_sc_hd__mux2_1 _4997_ (.A0(_2484_),
    .A1(_2485_),
    .S(net416),
    .X(_2486_));
 sky130_fd_sc_hd__mux4_1 _4998_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ),
    .S0(net434),
    .S1(net424),
    .X(_2487_));
 sky130_fd_sc_hd__mux4_1 _4999_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ),
    .S0(net431),
    .S1(net424),
    .X(_2488_));
 sky130_fd_sc_hd__mux2_1 _5000_ (.A0(_2488_),
    .A1(_2487_),
    .S(net414),
    .X(_2489_));
 sky130_fd_sc_hd__mux2_1 _5001_ (.A0(_2489_),
    .A1(_2486_),
    .S(net409),
    .X(_0058_));
 sky130_fd_sc_hd__mux4_1 _5002_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ),
    .S0(net433),
    .S1(net422),
    .X(_2490_));
 sky130_fd_sc_hd__mux4_1 _5003_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ),
    .S0(net436),
    .S1(net422),
    .X(_2491_));
 sky130_fd_sc_hd__mux2_1 _5004_ (.A0(_2490_),
    .A1(_2491_),
    .S(net414),
    .X(_2492_));
 sky130_fd_sc_hd__mux4_1 _5005_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ),
    .S0(net433),
    .S1(net422),
    .X(_2493_));
 sky130_fd_sc_hd__mux4_1 _5006_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ),
    .S0(net433),
    .S1(net422),
    .X(_2494_));
 sky130_fd_sc_hd__mux2_1 _5007_ (.A0(_2494_),
    .A1(_2493_),
    .S(net414),
    .X(_2495_));
 sky130_fd_sc_hd__mux2_1 _5008_ (.A0(_2495_),
    .A1(_2492_),
    .S(net409),
    .X(_0059_));
 sky130_fd_sc_hd__mux4_1 _5009_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ),
    .S0(net431),
    .S1(net421),
    .X(_2496_));
 sky130_fd_sc_hd__mux4_1 _5010_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ),
    .S0(net431),
    .S1(net421),
    .X(_2497_));
 sky130_fd_sc_hd__mux2_1 _5011_ (.A0(_2496_),
    .A1(_2497_),
    .S(net416),
    .X(_2498_));
 sky130_fd_sc_hd__mux4_1 _5012_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ),
    .S0(net431),
    .S1(net421),
    .X(_2499_));
 sky130_fd_sc_hd__mux4_1 _5013_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ),
    .S0(net431),
    .S1(net421),
    .X(_2500_));
 sky130_fd_sc_hd__mux2_1 _5014_ (.A0(_2500_),
    .A1(_2499_),
    .S(net416),
    .X(_2501_));
 sky130_fd_sc_hd__mux2_1 _5015_ (.A0(_2501_),
    .A1(_2498_),
    .S(net409),
    .X(_0060_));
 sky130_fd_sc_hd__mux4_1 _5016_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ),
    .S0(net427),
    .S1(net417),
    .X(_2502_));
 sky130_fd_sc_hd__mux4_1 _5017_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ),
    .S0(net428),
    .S1(net418),
    .X(_2503_));
 sky130_fd_sc_hd__mux2_1 _5018_ (.A0(_2502_),
    .A1(_2503_),
    .S(net411),
    .X(_2504_));
 sky130_fd_sc_hd__mux4_1 _5019_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ),
    .S0(net428),
    .S1(net418),
    .X(_2505_));
 sky130_fd_sc_hd__mux4_1 _5020_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ),
    .S0(net428),
    .S1(net417),
    .X(_2506_));
 sky130_fd_sc_hd__mux2_1 _5021_ (.A0(_2506_),
    .A1(_2505_),
    .S(net411),
    .X(_2507_));
 sky130_fd_sc_hd__mux2_1 _5022_ (.A0(_2507_),
    .A1(_2504_),
    .S(net410),
    .X(_0061_));
 sky130_fd_sc_hd__mux4_1 _5023_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ),
    .S0(net428),
    .S1(net418),
    .X(_2508_));
 sky130_fd_sc_hd__mux4_1 _5024_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ),
    .S0(net428),
    .S1(net418),
    .X(_2509_));
 sky130_fd_sc_hd__mux2_1 _5025_ (.A0(_2508_),
    .A1(_2509_),
    .S(net411),
    .X(_2510_));
 sky130_fd_sc_hd__mux4_1 _5026_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .S1(net426),
    .X(_2511_));
 sky130_fd_sc_hd__mux4_1 _5027_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ),
    .S0(net430),
    .S1(net420),
    .X(_2512_));
 sky130_fd_sc_hd__mux2_1 _5028_ (.A0(_2512_),
    .A1(_2511_),
    .S(net413),
    .X(_2513_));
 sky130_fd_sc_hd__mux2_1 _5029_ (.A0(_2513_),
    .A1(_2510_),
    .S(net410),
    .X(_0062_));
 sky130_fd_sc_hd__mux4_1 _5030_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ),
    .S0(net432),
    .S1(net421),
    .X(_2514_));
 sky130_fd_sc_hd__mux4_1 _5031_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ),
    .S0(net432),
    .S1(net421),
    .X(_2515_));
 sky130_fd_sc_hd__mux2_1 _5032_ (.A0(_2514_),
    .A1(_2515_),
    .S(net416),
    .X(_2516_));
 sky130_fd_sc_hd__mux4_1 _5033_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ),
    .S0(net431),
    .S1(net421),
    .X(_2517_));
 sky130_fd_sc_hd__mux4_1 _5034_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ),
    .S0(net431),
    .S1(net421),
    .X(_2518_));
 sky130_fd_sc_hd__mux2_1 _5035_ (.A0(_2518_),
    .A1(_2517_),
    .S(net416),
    .X(_2519_));
 sky130_fd_sc_hd__mux2_1 _5036_ (.A0(_2519_),
    .A1(_2516_),
    .S(net409),
    .X(_0063_));
 sky130_fd_sc_hd__mux4_1 _5037_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .S1(net426),
    .X(_2520_));
 sky130_fd_sc_hd__mux4_1 _5038_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .S1(net426),
    .X(_2521_));
 sky130_fd_sc_hd__mux2_1 _5039_ (.A0(_2520_),
    .A1(_2521_),
    .S(net413),
    .X(_2522_));
 sky130_fd_sc_hd__mux4_1 _5040_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ),
    .S0(net430),
    .S1(net420),
    .X(_2523_));
 sky130_fd_sc_hd__mux4_1 _5041_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .S1(net420),
    .X(_2524_));
 sky130_fd_sc_hd__mux2_1 _5042_ (.A0(_2524_),
    .A1(_2523_),
    .S(net413),
    .X(_2525_));
 sky130_fd_sc_hd__mux2_1 _5043_ (.A0(_2525_),
    .A1(_2522_),
    .S(net410),
    .X(_0033_));
 sky130_fd_sc_hd__mux4_1 _5044_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ),
    .S0(net428),
    .S1(net418),
    .X(_2526_));
 sky130_fd_sc_hd__mux4_1 _5045_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ),
    .S0(net427),
    .S1(net418),
    .X(_2527_));
 sky130_fd_sc_hd__mux2_1 _5046_ (.A0(_2526_),
    .A1(_2527_),
    .S(net411),
    .X(_2528_));
 sky130_fd_sc_hd__mux4_1 _5047_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ),
    .S0(net428),
    .S1(net418),
    .X(_2529_));
 sky130_fd_sc_hd__mux4_1 _5048_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ),
    .S0(net428),
    .S1(net418),
    .X(_2530_));
 sky130_fd_sc_hd__mux2_1 _5049_ (.A0(_2530_),
    .A1(_2529_),
    .S(net411),
    .X(_2531_));
 sky130_fd_sc_hd__mux2_1 _5050_ (.A0(_2531_),
    .A1(_2528_),
    .S(net410),
    .X(_0034_));
 sky130_fd_sc_hd__mux4_1 _5051_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ),
    .S0(net431),
    .S1(net421),
    .X(_2532_));
 sky130_fd_sc_hd__mux4_1 _5052_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ),
    .S0(net431),
    .S1(net424),
    .X(_2533_));
 sky130_fd_sc_hd__mux2_1 _5053_ (.A0(_2532_),
    .A1(_2533_),
    .S(net414),
    .X(_2534_));
 sky130_fd_sc_hd__mux4_1 _5054_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ),
    .S0(net431),
    .S1(net426),
    .X(_2535_));
 sky130_fd_sc_hd__mux4_1 _5055_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ),
    .S0(net431),
    .S1(net426),
    .X(_2536_));
 sky130_fd_sc_hd__mux2_1 _5056_ (.A0(_2536_),
    .A1(_2535_),
    .S(net416),
    .X(_2537_));
 sky130_fd_sc_hd__mux2_1 _5057_ (.A0(_2537_),
    .A1(_2534_),
    .S(net409),
    .X(_0035_));
 sky130_fd_sc_hd__mux4_1 _5058_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ),
    .S0(net431),
    .S1(net421),
    .X(_2538_));
 sky130_fd_sc_hd__mux4_1 _5059_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ),
    .S0(net434),
    .S1(net424),
    .X(_2539_));
 sky130_fd_sc_hd__mux2_1 _5060_ (.A0(_2538_),
    .A1(_2539_),
    .S(net414),
    .X(_2540_));
 sky130_fd_sc_hd__mux4_1 _5061_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ),
    .S0(net434),
    .S1(net424),
    .X(_2541_));
 sky130_fd_sc_hd__mux4_1 _5062_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ),
    .S0(net431),
    .S1(net421),
    .X(_2542_));
 sky130_fd_sc_hd__mux2_1 _5063_ (.A0(_2542_),
    .A1(_2541_),
    .S(net415),
    .X(_2543_));
 sky130_fd_sc_hd__mux2_1 _5064_ (.A0(_2543_),
    .A1(_2540_),
    .S(net409),
    .X(_0036_));
 sky130_fd_sc_hd__mux4_1 _5065_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ),
    .S0(net433),
    .S1(net425),
    .X(_2544_));
 sky130_fd_sc_hd__mux4_1 _5066_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ),
    .S0(net436),
    .S1(net425),
    .X(_2545_));
 sky130_fd_sc_hd__mux2_1 _5067_ (.A0(_2544_),
    .A1(_2545_),
    .S(net414),
    .X(_2546_));
 sky130_fd_sc_hd__mux4_1 _5068_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ),
    .S0(net433),
    .S1(net425),
    .X(_2547_));
 sky130_fd_sc_hd__mux4_1 _5069_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ),
    .S0(net433),
    .S1(net425),
    .X(_2548_));
 sky130_fd_sc_hd__mux2_1 _5070_ (.A0(_2548_),
    .A1(_2547_),
    .S(net414),
    .X(_2549_));
 sky130_fd_sc_hd__mux2_1 _5071_ (.A0(_2549_),
    .A1(_2546_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .X(_0037_));
 sky130_fd_sc_hd__mux4_1 _5072_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ),
    .S0(net432),
    .S1(net422),
    .X(_2550_));
 sky130_fd_sc_hd__mux4_1 _5073_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ),
    .S0(net433),
    .S1(net422),
    .X(_2551_));
 sky130_fd_sc_hd__mux2_1 _5074_ (.A0(_2550_),
    .A1(_2551_),
    .S(net414),
    .X(_2552_));
 sky130_fd_sc_hd__mux4_1 _5075_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ),
    .S0(net433),
    .S1(net422),
    .X(_2553_));
 sky130_fd_sc_hd__mux4_1 _5076_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ),
    .S0(net432),
    .S1(net422),
    .X(_2554_));
 sky130_fd_sc_hd__mux2_1 _5077_ (.A0(_2554_),
    .A1(_2553_),
    .S(net414),
    .X(_2555_));
 sky130_fd_sc_hd__mux2_1 _5078_ (.A0(_2555_),
    .A1(_2552_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .X(_0038_));
 sky130_fd_sc_hd__mux4_1 _5079_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ),
    .S0(net430),
    .S1(net420),
    .X(_2556_));
 sky130_fd_sc_hd__mux4_1 _5080_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ),
    .S0(net430),
    .S1(net420),
    .X(_2557_));
 sky130_fd_sc_hd__mux2_1 _5081_ (.A0(_2556_),
    .A1(_2557_),
    .S(net413),
    .X(_2558_));
 sky130_fd_sc_hd__mux4_1 _5082_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ),
    .S0(net430),
    .S1(net420),
    .X(_2559_));
 sky130_fd_sc_hd__mux4_1 _5083_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ),
    .S0(net430),
    .S1(net420),
    .X(_2560_));
 sky130_fd_sc_hd__mux2_1 _5084_ (.A0(_2560_),
    .A1(_2559_),
    .S(net413),
    .X(_2561_));
 sky130_fd_sc_hd__mux2_1 _5085_ (.A0(_2561_),
    .A1(_2558_),
    .S(net410),
    .X(_0039_));
 sky130_fd_sc_hd__mux4_1 _5086_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ),
    .S0(net431),
    .S1(net421),
    .X(_2562_));
 sky130_fd_sc_hd__mux4_1 _5087_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ),
    .S0(net431),
    .S1(net421),
    .X(_2563_));
 sky130_fd_sc_hd__mux2_1 _5088_ (.A0(_2562_),
    .A1(_2563_),
    .S(net416),
    .X(_2564_));
 sky130_fd_sc_hd__mux4_1 _5089_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ),
    .S0(net431),
    .S1(net421),
    .X(_2565_));
 sky130_fd_sc_hd__mux4_1 _5090_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ),
    .S0(net430),
    .S1(net420),
    .X(_2566_));
 sky130_fd_sc_hd__mux2_1 _5091_ (.A0(_2566_),
    .A1(_2565_),
    .S(net416),
    .X(_2567_));
 sky130_fd_sc_hd__mux2_1 _5092_ (.A0(_2567_),
    .A1(_2564_),
    .S(net409),
    .X(_0040_));
 sky130_fd_sc_hd__mux4_1 _5093_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ),
    .S0(net436),
    .S1(net422),
    .X(_2568_));
 sky130_fd_sc_hd__mux4_1 _5094_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ),
    .S0(net436),
    .S1(net422),
    .X(_2569_));
 sky130_fd_sc_hd__mux2_1 _5095_ (.A0(_2568_),
    .A1(_2569_),
    .S(net414),
    .X(_2570_));
 sky130_fd_sc_hd__mux4_1 _5096_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ),
    .S0(net436),
    .S1(net422),
    .X(_2571_));
 sky130_fd_sc_hd__mux4_1 _5097_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ),
    .S0(net433),
    .S1(net425),
    .X(_2572_));
 sky130_fd_sc_hd__mux2_1 _5098_ (.A0(_2572_),
    .A1(_2571_),
    .S(net414),
    .X(_2573_));
 sky130_fd_sc_hd__mux2_1 _5099_ (.A0(_2573_),
    .A1(_2570_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .X(_0041_));
 sky130_fd_sc_hd__mux4_1 _5100_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ),
    .S0(net433),
    .S1(net422),
    .X(_2574_));
 sky130_fd_sc_hd__mux4_1 _5101_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ),
    .S0(net433),
    .S1(net422),
    .X(_2575_));
 sky130_fd_sc_hd__mux2_1 _5102_ (.A0(_2574_),
    .A1(_2575_),
    .S(net414),
    .X(_2576_));
 sky130_fd_sc_hd__mux4_1 _5103_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ),
    .S0(net432),
    .S1(net422),
    .X(_2577_));
 sky130_fd_sc_hd__mux4_1 _5104_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ),
    .S0(net433),
    .S1(net422),
    .X(_2578_));
 sky130_fd_sc_hd__mux2_1 _5105_ (.A0(_2578_),
    .A1(_2577_),
    .S(net414),
    .X(_2579_));
 sky130_fd_sc_hd__mux2_1 _5106_ (.A0(_2579_),
    .A1(_2576_),
    .S(net409),
    .X(_0042_));
 sky130_fd_sc_hd__mux4_1 _5107_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ),
    .S0(net429),
    .S1(net419),
    .X(_2580_));
 sky130_fd_sc_hd__mux4_1 _5108_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ),
    .S0(net429),
    .S1(net419),
    .X(_2581_));
 sky130_fd_sc_hd__mux2_1 _5109_ (.A0(_2580_),
    .A1(_2581_),
    .S(net412),
    .X(_2582_));
 sky130_fd_sc_hd__mux4_1 _5110_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ),
    .S0(net429),
    .S1(net419),
    .X(_2583_));
 sky130_fd_sc_hd__mux4_1 _5111_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ),
    .S0(net429),
    .S1(net419),
    .X(_2584_));
 sky130_fd_sc_hd__mux2_1 _5112_ (.A0(_2584_),
    .A1(_2583_),
    .S(net412),
    .X(_2585_));
 sky130_fd_sc_hd__mux2_1 _5113_ (.A0(_2585_),
    .A1(_2582_),
    .S(net410),
    .X(_0044_));
 sky130_fd_sc_hd__mux4_1 _5114_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ),
    .S0(net429),
    .S1(net419),
    .X(_2586_));
 sky130_fd_sc_hd__mux4_1 _5115_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ),
    .S0(net429),
    .S1(net419),
    .X(_2587_));
 sky130_fd_sc_hd__mux2_1 _5116_ (.A0(_2586_),
    .A1(_2587_),
    .S(net412),
    .X(_2588_));
 sky130_fd_sc_hd__mux4_1 _5117_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ),
    .S0(net429),
    .S1(net419),
    .X(_2589_));
 sky130_fd_sc_hd__mux4_1 _5118_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ),
    .S0(net429),
    .S1(net419),
    .X(_2590_));
 sky130_fd_sc_hd__mux2_1 _5119_ (.A0(_2590_),
    .A1(_2589_),
    .S(net412),
    .X(_2591_));
 sky130_fd_sc_hd__mux2_1 _5120_ (.A0(_2591_),
    .A1(_2588_),
    .S(net410),
    .X(_0045_));
 sky130_fd_sc_hd__mux4_1 _5121_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ),
    .S0(net434),
    .S1(net424),
    .X(_2592_));
 sky130_fd_sc_hd__mux4_1 _5122_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ),
    .S0(net434),
    .S1(net424),
    .X(_2593_));
 sky130_fd_sc_hd__mux2_1 _5123_ (.A0(_2592_),
    .A1(_2593_),
    .S(net415),
    .X(_2594_));
 sky130_fd_sc_hd__mux4_1 _5124_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ),
    .S0(net434),
    .S1(net424),
    .X(_2595_));
 sky130_fd_sc_hd__mux4_1 _5125_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ),
    .S0(net434),
    .S1(net424),
    .X(_2596_));
 sky130_fd_sc_hd__mux2_1 _5126_ (.A0(_2596_),
    .A1(_2595_),
    .S(net415),
    .X(_2597_));
 sky130_fd_sc_hd__mux2_1 _5127_ (.A0(_2597_),
    .A1(_2594_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .X(_0046_));
 sky130_fd_sc_hd__mux4_1 _5128_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ),
    .S0(net429),
    .S1(net419),
    .X(_2598_));
 sky130_fd_sc_hd__mux4_1 _5129_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ),
    .S0(net427),
    .S1(net418),
    .X(_2599_));
 sky130_fd_sc_hd__mux2_1 _5130_ (.A0(_2598_),
    .A1(_2599_),
    .S(net411),
    .X(_2600_));
 sky130_fd_sc_hd__mux4_1 _5131_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ),
    .S0(net429),
    .S1(net419),
    .X(_2601_));
 sky130_fd_sc_hd__mux4_1 _5132_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ),
    .S0(net429),
    .S1(net419),
    .X(_2602_));
 sky130_fd_sc_hd__mux2_1 _5133_ (.A0(_2602_),
    .A1(_2601_),
    .S(net411),
    .X(_2603_));
 sky130_fd_sc_hd__mux2_1 _5134_ (.A0(_2603_),
    .A1(_2600_),
    .S(net410),
    .X(_0047_));
 sky130_fd_sc_hd__mux4_1 _5135_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ),
    .S0(net434),
    .S1(net424),
    .X(_2604_));
 sky130_fd_sc_hd__mux4_1 _5136_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ),
    .S0(net434),
    .S1(net424),
    .X(_2605_));
 sky130_fd_sc_hd__mux2_1 _5137_ (.A0(_2604_),
    .A1(_2605_),
    .S(net415),
    .X(_2606_));
 sky130_fd_sc_hd__mux4_1 _5138_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ),
    .S0(net434),
    .S1(net424),
    .X(_2607_));
 sky130_fd_sc_hd__mux4_1 _5139_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ),
    .S0(net434),
    .S1(net424),
    .X(_2608_));
 sky130_fd_sc_hd__mux2_1 _5140_ (.A0(_2608_),
    .A1(_2607_),
    .S(net415),
    .X(_2609_));
 sky130_fd_sc_hd__mux2_1 _5141_ (.A0(_2609_),
    .A1(_2606_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .X(_0048_));
 sky130_fd_sc_hd__mux4_1 _5142_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ),
    .S0(net427),
    .S1(net417),
    .X(_2610_));
 sky130_fd_sc_hd__mux4_1 _5143_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ),
    .S0(net427),
    .S1(net417),
    .X(_2611_));
 sky130_fd_sc_hd__mux2_1 _5144_ (.A0(_2610_),
    .A1(_2611_),
    .S(net411),
    .X(_2612_));
 sky130_fd_sc_hd__mux4_1 _5145_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ),
    .S0(net427),
    .S1(net417),
    .X(_2613_));
 sky130_fd_sc_hd__mux4_1 _5146_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ),
    .S0(net428),
    .S1(net417),
    .X(_2614_));
 sky130_fd_sc_hd__mux2_1 _5147_ (.A0(_2614_),
    .A1(_2613_),
    .S(net411),
    .X(_2615_));
 sky130_fd_sc_hd__mux2_1 _5148_ (.A0(_2615_),
    .A1(_2612_),
    .S(net410),
    .X(_0049_));
 sky130_fd_sc_hd__mux4_1 _5149_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ),
    .S0(net429),
    .S1(net419),
    .X(_2616_));
 sky130_fd_sc_hd__mux4_1 _5150_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ),
    .S0(net429),
    .S1(net419),
    .X(_2617_));
 sky130_fd_sc_hd__mux2_1 _5151_ (.A0(_2616_),
    .A1(_2617_),
    .S(net412),
    .X(_2618_));
 sky130_fd_sc_hd__mux4_1 _5152_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ),
    .S0(net429),
    .S1(net419),
    .X(_2619_));
 sky130_fd_sc_hd__mux4_1 _5153_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ),
    .S0(net429),
    .S1(net419),
    .X(_2620_));
 sky130_fd_sc_hd__mux2_1 _5154_ (.A0(_2620_),
    .A1(_2619_),
    .S(net412),
    .X(_2621_));
 sky130_fd_sc_hd__mux2_1 _5155_ (.A0(_2621_),
    .A1(_2618_),
    .S(net410),
    .X(_0050_));
 sky130_fd_sc_hd__mux4_1 _5156_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ),
    .S0(net430),
    .S1(net421),
    .X(_2622_));
 sky130_fd_sc_hd__mux4_1 _5157_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ),
    .S0(net430),
    .S1(net420),
    .X(_2623_));
 sky130_fd_sc_hd__mux2_1 _5158_ (.A0(_2622_),
    .A1(_2623_),
    .S(net413),
    .X(_2624_));
 sky130_fd_sc_hd__mux4_1 _5159_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ),
    .S0(net430),
    .S1(net420),
    .X(_2625_));
 sky130_fd_sc_hd__mux4_1 _5160_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ),
    .S0(net430),
    .S1(net421),
    .X(_2626_));
 sky130_fd_sc_hd__mux2_1 _5161_ (.A0(_2626_),
    .A1(_2625_),
    .S(net413),
    .X(_2627_));
 sky130_fd_sc_hd__mux2_1 _5162_ (.A0(_2627_),
    .A1(_2624_),
    .S(net410),
    .X(_0051_));
 sky130_fd_sc_hd__mux4_1 _5163_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ),
    .S0(net427),
    .S1(net417),
    .X(_2628_));
 sky130_fd_sc_hd__mux4_1 _5164_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ),
    .S0(net427),
    .S1(net417),
    .X(_2629_));
 sky130_fd_sc_hd__mux2_1 _5165_ (.A0(_2628_),
    .A1(_2629_),
    .S(net411),
    .X(_2630_));
 sky130_fd_sc_hd__mux4_1 _5166_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ),
    .S0(net427),
    .S1(net417),
    .X(_2631_));
 sky130_fd_sc_hd__mux4_1 _5167_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ),
    .S0(net427),
    .S1(net417),
    .X(_2632_));
 sky130_fd_sc_hd__mux2_1 _5168_ (.A0(_2632_),
    .A1(_2631_),
    .S(net411),
    .X(_2633_));
 sky130_fd_sc_hd__mux2_1 _5169_ (.A0(_2633_),
    .A1(_2630_),
    .S(net410),
    .X(_0052_));
 sky130_fd_sc_hd__mux4_1 _5170_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ),
    .S0(net428),
    .S1(net418),
    .X(_2634_));
 sky130_fd_sc_hd__mux4_1 _5171_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ),
    .S0(net428),
    .S1(net418),
    .X(_2635_));
 sky130_fd_sc_hd__mux2_1 _5172_ (.A0(_2634_),
    .A1(_2635_),
    .S(net411),
    .X(_2636_));
 sky130_fd_sc_hd__mux4_1 _5173_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ),
    .S0(net427),
    .S1(net417),
    .X(_2637_));
 sky130_fd_sc_hd__mux4_1 _5174_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ),
    .S0(net427),
    .S1(net417),
    .X(_2638_));
 sky130_fd_sc_hd__mux2_1 _5175_ (.A0(_2638_),
    .A1(_2637_),
    .S(net411),
    .X(_2639_));
 sky130_fd_sc_hd__mux2_1 _5176_ (.A0(_2639_),
    .A1(_2636_),
    .S(net410),
    .X(_0053_));
 sky130_fd_sc_hd__mux4_1 _5177_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ),
    .S0(net427),
    .S1(net417),
    .X(_2640_));
 sky130_fd_sc_hd__mux4_1 _5178_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ),
    .S0(net427),
    .S1(net417),
    .X(_2641_));
 sky130_fd_sc_hd__mux2_1 _5179_ (.A0(_2640_),
    .A1(_2641_),
    .S(net411),
    .X(_2642_));
 sky130_fd_sc_hd__mux4_1 _5180_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ),
    .S0(net427),
    .S1(net417),
    .X(_2643_));
 sky130_fd_sc_hd__mux4_1 _5181_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ),
    .S0(net427),
    .S1(net417),
    .X(_2644_));
 sky130_fd_sc_hd__mux2_1 _5182_ (.A0(_2644_),
    .A1(_2643_),
    .S(net411),
    .X(_2645_));
 sky130_fd_sc_hd__mux2_1 _5183_ (.A0(_2645_),
    .A1(_2642_),
    .S(net410),
    .X(_0055_));
 sky130_fd_sc_hd__mux4_1 _5184_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ),
    .S0(net430),
    .S1(net419),
    .X(_2646_));
 sky130_fd_sc_hd__mux4_1 _5185_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ),
    .S0(net430),
    .S1(net420),
    .X(_2647_));
 sky130_fd_sc_hd__mux2_1 _5186_ (.A0(_2646_),
    .A1(_2647_),
    .S(net412),
    .X(_2648_));
 sky130_fd_sc_hd__mux4_1 _5187_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ),
    .S0(net429),
    .S1(net420),
    .X(_2649_));
 sky130_fd_sc_hd__mux4_1 _5188_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ),
    .S0(net430),
    .S1(net420),
    .X(_2650_));
 sky130_fd_sc_hd__mux2_1 _5189_ (.A0(_2650_),
    .A1(_2649_),
    .S(net412),
    .X(_2651_));
 sky130_fd_sc_hd__mux2_1 _5190_ (.A0(_2651_),
    .A1(_2648_),
    .S(net410),
    .X(_0056_));
 sky130_fd_sc_hd__and2_1 _5191_ (.A(net452),
    .B(net789),
    .X(_0290_));
 sky130_fd_sc_hd__and2_1 _5192_ (.A(net456),
    .B(net715),
    .X(_0291_));
 sky130_fd_sc_hd__and2_1 _5193_ (.A(net466),
    .B(net182),
    .X(_2652_));
 sky130_fd_sc_hd__mux2_1 _5194_ (.A0(net2131),
    .A1(net801),
    .S(net301),
    .X(_2653_));
 sky130_fd_sc_hd__or3b_1 _5195_ (.A(net480),
    .B(_2653_),
    .C_N(net183),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _5196_ (.A(net946),
    .B(net288),
    .X(_2654_));
 sky130_fd_sc_hd__o211a_1 _5197_ (.A1(net2052),
    .A2(net301),
    .B1(net168),
    .C1(_2654_),
    .X(_0323_));
 sky130_fd_sc_hd__or2_1 _5198_ (.A(net992),
    .B(net288),
    .X(_2655_));
 sky130_fd_sc_hd__o211a_1 _5199_ (.A1(net2013),
    .A2(net301),
    .B1(net168),
    .C1(_2655_),
    .X(_0324_));
 sky130_fd_sc_hd__or2_1 _5200_ (.A(net894),
    .B(net282),
    .X(_2656_));
 sky130_fd_sc_hd__o211a_1 _5201_ (.A1(net2005),
    .A2(net299),
    .B1(net167),
    .C1(_2656_),
    .X(_0325_));
 sky130_fd_sc_hd__or2_1 _5202_ (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ),
    .B(net282),
    .X(_2657_));
 sky130_fd_sc_hd__o211a_1 _5203_ (.A1(net1982),
    .A2(net296),
    .B1(net166),
    .C1(_2657_),
    .X(_0326_));
 sky130_fd_sc_hd__or2_1 _5204_ (.A(net944),
    .B(net277),
    .X(_2658_));
 sky130_fd_sc_hd__o211a_1 _5205_ (.A1(net1969),
    .A2(net296),
    .B1(net166),
    .C1(_2658_),
    .X(_0327_));
 sky130_fd_sc_hd__or2_1 _5206_ (.A(net896),
    .B(net282),
    .X(_2659_));
 sky130_fd_sc_hd__o211a_1 _5207_ (.A1(net2033),
    .A2(net297),
    .B1(net166),
    .C1(_2659_),
    .X(_0328_));
 sky130_fd_sc_hd__or2_1 _5208_ (.A(net932),
    .B(net282),
    .X(_2660_));
 sky130_fd_sc_hd__o211a_1 _5209_ (.A1(net2001),
    .A2(net299),
    .B1(net167),
    .C1(_2660_),
    .X(_0329_));
 sky130_fd_sc_hd__or2_1 _5210_ (.A(net902),
    .B(net279),
    .X(_2661_));
 sky130_fd_sc_hd__o211a_1 _5211_ (.A1(net2038),
    .A2(net297),
    .B1(net166),
    .C1(_2661_),
    .X(_0330_));
 sky130_fd_sc_hd__or2_1 _5212_ (.A(net868),
    .B(net279),
    .X(_2662_));
 sky130_fd_sc_hd__o211a_1 _5213_ (.A1(net1996),
    .A2(net297),
    .B1(net166),
    .C1(_2662_),
    .X(_0331_));
 sky130_fd_sc_hd__or2_1 _5214_ (.A(net922),
    .B(net277),
    .X(_2663_));
 sky130_fd_sc_hd__o211a_1 _5215_ (.A1(net1949),
    .A2(net296),
    .B1(net166),
    .C1(_2663_),
    .X(_0332_));
 sky130_fd_sc_hd__or2_1 _5216_ (.A(net974),
    .B(net283),
    .X(_2664_));
 sky130_fd_sc_hd__o211a_1 _5217_ (.A1(net2048),
    .A2(net299),
    .B1(net167),
    .C1(_2664_),
    .X(_0333_));
 sky130_fd_sc_hd__or2_1 _5218_ (.A(net960),
    .B(net283),
    .X(_2665_));
 sky130_fd_sc_hd__o211a_1 _5219_ (.A1(net2028),
    .A2(net299),
    .B1(net167),
    .C1(_2665_),
    .X(_0334_));
 sky130_fd_sc_hd__or2_1 _5220_ (.A(net964),
    .B(net285),
    .X(_2666_));
 sky130_fd_sc_hd__o211a_1 _5221_ (.A1(net2017),
    .A2(net300),
    .B1(net169),
    .C1(_2666_),
    .X(_0335_));
 sky130_fd_sc_hd__or2_1 _5222_ (.A(net2086),
    .B(net285),
    .X(_2667_));
 sky130_fd_sc_hd__o211a_1 _5223_ (.A1(net2042),
    .A2(net299),
    .B1(net167),
    .C1(_2667_),
    .X(_0336_));
 sky130_fd_sc_hd__or2_1 _5224_ (.A(net1331),
    .B(net285),
    .X(_2668_));
 sky130_fd_sc_hd__o211a_1 _5225_ (.A1(net2079),
    .A2(net300),
    .B1(net167),
    .C1(_2668_),
    .X(_0337_));
 sky130_fd_sc_hd__or2_1 _5226_ (.A(net713),
    .B(net289),
    .X(_2669_));
 sky130_fd_sc_hd__o211a_1 _5227_ (.A1(net2030),
    .A2(net301),
    .B1(net168),
    .C1(_2669_),
    .X(_0338_));
 sky130_fd_sc_hd__or2_1 _5228_ (.A(net1315),
    .B(net285),
    .X(_2670_));
 sky130_fd_sc_hd__o211a_1 _5229_ (.A1(net1333),
    .A2(net300),
    .B1(net167),
    .C1(_2670_),
    .X(_0339_));
 sky130_fd_sc_hd__or2_1 _5230_ (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[20] ),
    .B(net292),
    .X(_2671_));
 sky130_fd_sc_hd__o211a_1 _5231_ (.A1(net735),
    .A2(net302),
    .B1(net169),
    .C1(_2671_),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _5232_ (.A(net1132),
    .B(net276),
    .X(_2672_));
 sky130_fd_sc_hd__o211a_1 _5233_ (.A1(net1828),
    .A2(net294),
    .B1(net164),
    .C1(_2672_),
    .X(_0341_));
 sky130_fd_sc_hd__or2_1 _5234_ (.A(net942),
    .B(net276),
    .X(_2673_));
 sky130_fd_sc_hd__o211a_1 _5235_ (.A1(net2016),
    .A2(net298),
    .B1(net165),
    .C1(_2673_),
    .X(_0342_));
 sky130_fd_sc_hd__or2_1 _5236_ (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[23] ),
    .B(net276),
    .X(_2674_));
 sky130_fd_sc_hd__o211a_1 _5237_ (.A1(net661),
    .A2(net294),
    .B1(net164),
    .C1(_2674_),
    .X(_0343_));
 sky130_fd_sc_hd__or2_1 _5238_ (.A(net870),
    .B(net280),
    .X(_2675_));
 sky130_fd_sc_hd__o211a_1 _5239_ (.A1(net2072),
    .A2(net298),
    .B1(net170),
    .C1(_2675_),
    .X(_0344_));
 sky130_fd_sc_hd__or2_1 _5240_ (.A(net1004),
    .B(net274),
    .X(_2676_));
 sky130_fd_sc_hd__o211a_1 _5241_ (.A1(net2098),
    .A2(net293),
    .B1(net164),
    .C1(_2676_),
    .X(_0345_));
 sky130_fd_sc_hd__or2_1 _5242_ (.A(net1076),
    .B(net275),
    .X(_2677_));
 sky130_fd_sc_hd__o211a_1 _5243_ (.A1(net2087),
    .A2(net293),
    .B1(net164),
    .C1(_2677_),
    .X(_0346_));
 sky130_fd_sc_hd__or2_1 _5244_ (.A(net1108),
    .B(net276),
    .X(_2678_));
 sky130_fd_sc_hd__o211a_1 _5245_ (.A1(net2060),
    .A2(net294),
    .B1(net164),
    .C1(_2678_),
    .X(_0347_));
 sky130_fd_sc_hd__or2_1 _5246_ (.A(net671),
    .B(net272),
    .X(_2679_));
 sky130_fd_sc_hd__o211a_1 _5247_ (.A1(net2043),
    .A2(net295),
    .B1(net165),
    .C1(_2679_),
    .X(_0348_));
 sky130_fd_sc_hd__or2_1 _5248_ (.A(net1028),
    .B(net273),
    .X(_2680_));
 sky130_fd_sc_hd__o211a_1 _5249_ (.A1(net2049),
    .A2(net295),
    .B1(net165),
    .C1(_2680_),
    .X(_0349_));
 sky130_fd_sc_hd__or2_1 _5250_ (.A(net1810),
    .B(net273),
    .X(_2681_));
 sky130_fd_sc_hd__o211a_1 _5251_ (.A1(net2070),
    .A2(net295),
    .B1(net165),
    .C1(_2681_),
    .X(_0350_));
 sky130_fd_sc_hd__or2_1 _5252_ (.A(net1020),
    .B(net280),
    .X(_2682_));
 sky130_fd_sc_hd__o211a_1 _5253_ (.A1(net1850),
    .A2(net294),
    .B1(net164),
    .C1(_2682_),
    .X(_0351_));
 sky130_fd_sc_hd__nand2_1 _5254_ (.A(_1408_),
    .B(net296),
    .Y(_2683_));
 sky130_fd_sc_hd__o211a_1 _5255_ (.A1(net21),
    .A2(net296),
    .B1(net166),
    .C1(_2683_),
    .X(_0352_));
 sky130_fd_sc_hd__or2_1 _5256_ (.A(net2058),
    .B(net277),
    .X(_2684_));
 sky130_fd_sc_hd__o211a_1 _5257_ (.A1(net24),
    .A2(net296),
    .B1(net166),
    .C1(_2684_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _5258_ (.A0(net25),
    .A1(net2203),
    .S(net296),
    .X(_2685_));
 sky130_fd_sc_hd__or3b_1 _5259_ (.A(net476),
    .B(_2685_),
    .C_N(net176),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _5260_ (.A0(net26),
    .A1(net2197),
    .S(net296),
    .X(_2686_));
 sky130_fd_sc_hd__or3b_1 _5261_ (.A(net476),
    .B(_2686_),
    .C_N(net176),
    .X(_0355_));
 sky130_fd_sc_hd__nand2_1 _5262_ (.A(_1407_),
    .B(net296),
    .Y(_2687_));
 sky130_fd_sc_hd__o211a_1 _5263_ (.A1(net27),
    .A2(net296),
    .B1(net166),
    .C1(_2687_),
    .X(_0356_));
 sky130_fd_sc_hd__or2_1 _5264_ (.A(net2128),
    .B(net290),
    .X(_2688_));
 sky130_fd_sc_hd__o211a_1 _5265_ (.A1(net28),
    .A2(net301),
    .B1(net168),
    .C1(_2688_),
    .X(_0357_));
 sky130_fd_sc_hd__or2_1 _5266_ (.A(net2204),
    .B(net282),
    .X(_2689_));
 sky130_fd_sc_hd__o211a_1 _5267_ (.A1(net29),
    .A2(net299),
    .B1(net167),
    .C1(_2689_),
    .X(_0358_));
 sky130_fd_sc_hd__or2_1 _5268_ (.A(net2103),
    .B(net291),
    .X(_2690_));
 sky130_fd_sc_hd__o211a_1 _5269_ (.A1(net30),
    .A2(net302),
    .B1(net168),
    .C1(_2690_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _5270_ (.A(net2134),
    .B(net290),
    .X(_2691_));
 sky130_fd_sc_hd__o211a_1 _5271_ (.A1(net1),
    .A2(net301),
    .B1(net168),
    .C1(_2691_),
    .X(_0360_));
 sky130_fd_sc_hd__or2_1 _5272_ (.A(net2199),
    .B(net277),
    .X(_2692_));
 sky130_fd_sc_hd__o211a_1 _5273_ (.A1(net2),
    .A2(net296),
    .B1(net166),
    .C1(_2692_),
    .X(_0361_));
 sky130_fd_sc_hd__or2_1 _5274_ (.A(net2010),
    .B(net280),
    .X(_2693_));
 sky130_fd_sc_hd__o211a_1 _5275_ (.A1(net3),
    .A2(net298),
    .B1(net170),
    .C1(_2693_),
    .X(_0362_));
 sky130_fd_sc_hd__or2_1 _5276_ (.A(net2092),
    .B(net290),
    .X(_2694_));
 sky130_fd_sc_hd__o211a_1 _5277_ (.A1(net4),
    .A2(net301),
    .B1(net168),
    .C1(_2694_),
    .X(_0363_));
 sky130_fd_sc_hd__or2_1 _5278_ (.A(net2055),
    .B(net289),
    .X(_2695_));
 sky130_fd_sc_hd__o211a_1 _5279_ (.A1(net5),
    .A2(net301),
    .B1(net168),
    .C1(_2695_),
    .X(_0364_));
 sky130_fd_sc_hd__or2_1 _5280_ (.A(net433),
    .B(net290),
    .X(_2696_));
 sky130_fd_sc_hd__o211a_1 _5281_ (.A1(net6),
    .A2(net301),
    .B1(net168),
    .C1(_2696_),
    .X(_0365_));
 sky130_fd_sc_hd__or2_1 _5282_ (.A(net420),
    .B(net280),
    .X(_2697_));
 sky130_fd_sc_hd__o211a_1 _5283_ (.A1(net7),
    .A2(net298),
    .B1(net170),
    .C1(_2697_),
    .X(_0366_));
 sky130_fd_sc_hd__or2_1 _5284_ (.A(net411),
    .B(net273),
    .X(_2698_));
 sky130_fd_sc_hd__o211a_1 _5285_ (.A1(net8),
    .A2(net293),
    .B1(net164),
    .C1(_2698_),
    .X(_0367_));
 sky130_fd_sc_hd__or2_1 _5286_ (.A(net410),
    .B(net272),
    .X(_2699_));
 sky130_fd_sc_hd__o211a_1 _5287_ (.A1(net9),
    .A2(net295),
    .B1(net165),
    .C1(_2699_),
    .X(_0368_));
 sky130_fd_sc_hd__or2_1 _5288_ (.A(net2105),
    .B(net291),
    .X(_2700_));
 sky130_fd_sc_hd__o211a_1 _5289_ (.A1(net10),
    .A2(net302),
    .B1(net168),
    .C1(_2700_),
    .X(_0369_));
 sky130_fd_sc_hd__or2_1 _5290_ (.A(net405),
    .B(net291),
    .X(_2701_));
 sky130_fd_sc_hd__o211a_1 _5291_ (.A1(net11),
    .A2(net302),
    .B1(net168),
    .C1(_2701_),
    .X(_0370_));
 sky130_fd_sc_hd__or2_1 _5292_ (.A(net392),
    .B(net276),
    .X(_2702_));
 sky130_fd_sc_hd__o211a_1 _5293_ (.A1(net12),
    .A2(net294),
    .B1(net164),
    .C1(_2702_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _5294_ (.A(net386),
    .B(net291),
    .X(_2703_));
 sky130_fd_sc_hd__o211a_1 _5295_ (.A1(net13),
    .A2(net302),
    .B1(net168),
    .C1(_2703_),
    .X(_0372_));
 sky130_fd_sc_hd__or2_1 _5296_ (.A(net381),
    .B(net275),
    .X(_2704_));
 sky130_fd_sc_hd__o211a_1 _5297_ (.A1(net14),
    .A2(net293),
    .B1(net164),
    .C1(_2704_),
    .X(_0373_));
 sky130_fd_sc_hd__or2_1 _5298_ (.A(net2172),
    .B(net292),
    .X(_2705_));
 sky130_fd_sc_hd__o211a_1 _5299_ (.A1(net15),
    .A2(net303),
    .B1(net169),
    .C1(_2705_),
    .X(_0374_));
 sky130_fd_sc_hd__or2_1 _5300_ (.A(net1292),
    .B(net279),
    .X(_2706_));
 sky130_fd_sc_hd__o211a_1 _5301_ (.A1(net16),
    .A2(net297),
    .B1(net166),
    .C1(_2706_),
    .X(_0375_));
 sky130_fd_sc_hd__or2_1 _5302_ (.A(net1997),
    .B(net272),
    .X(_2707_));
 sky130_fd_sc_hd__o211a_1 _5303_ (.A1(net17),
    .A2(net295),
    .B1(net165),
    .C1(_2707_),
    .X(_0376_));
 sky130_fd_sc_hd__or2_1 _5304_ (.A(net2214),
    .B(net291),
    .X(_2708_));
 sky130_fd_sc_hd__o211a_1 _5305_ (.A1(net18),
    .A2(net302),
    .B1(net169),
    .C1(_2708_),
    .X(_0377_));
 sky130_fd_sc_hd__or2_1 _5306_ (.A(net2007),
    .B(net272),
    .X(_2709_));
 sky130_fd_sc_hd__o211a_1 _5307_ (.A1(net19),
    .A2(net295),
    .B1(net165),
    .C1(_2709_),
    .X(_0378_));
 sky130_fd_sc_hd__or2_1 _5308_ (.A(net2138),
    .B(net290),
    .X(_2710_));
 sky130_fd_sc_hd__o211a_1 _5309_ (.A1(net20),
    .A2(net302),
    .B1(net168),
    .C1(_2710_),
    .X(_0379_));
 sky130_fd_sc_hd__or2_1 _5310_ (.A(net2190),
    .B(net275),
    .X(_2711_));
 sky130_fd_sc_hd__o211a_1 _5311_ (.A1(net22),
    .A2(net293),
    .B1(net164),
    .C1(_2711_),
    .X(_0380_));
 sky130_fd_sc_hd__or2_1 _5312_ (.A(net2019),
    .B(net279),
    .X(_2712_));
 sky130_fd_sc_hd__o211a_1 _5313_ (.A1(net23),
    .A2(net297),
    .B1(net166),
    .C1(_2712_),
    .X(_0381_));
 sky130_fd_sc_hd__or2_1 _5314_ (.A(net1357),
    .B(net288),
    .X(_2713_));
 sky130_fd_sc_hd__o211a_1 _5315_ (.A1(net2099),
    .A2(net301),
    .B1(net168),
    .C1(_2713_),
    .X(_0382_));
 sky130_fd_sc_hd__or2_1 _5316_ (.A(net627),
    .B(net290),
    .X(_2714_));
 sky130_fd_sc_hd__o211a_1 _5317_ (.A1(net2117),
    .A2(net301),
    .B1(net168),
    .C1(_2714_),
    .X(_0383_));
 sky130_fd_sc_hd__or2_1 _5318_ (.A(net882),
    .B(net284),
    .X(_2715_));
 sky130_fd_sc_hd__o211a_1 _5319_ (.A1(net2037),
    .A2(net299),
    .B1(net167),
    .C1(_2715_),
    .X(_0384_));
 sky130_fd_sc_hd__or2_1 _5320_ (.A(net978),
    .B(net282),
    .X(_2716_));
 sky130_fd_sc_hd__o211a_1 _5321_ (.A1(net2053),
    .A2(net299),
    .B1(net167),
    .C1(_2716_),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _5322_ (.A(net874),
    .B(net278),
    .X(_2717_));
 sky130_fd_sc_hd__o211a_1 _5323_ (.A1(net2026),
    .A2(net297),
    .B1(net166),
    .C1(_2717_),
    .X(_0386_));
 sky130_fd_sc_hd__or2_1 _5324_ (.A(net928),
    .B(net277),
    .X(_2718_));
 sky130_fd_sc_hd__o211a_1 _5325_ (.A1(net2063),
    .A2(net297),
    .B1(net166),
    .C1(_2718_),
    .X(_0387_));
 sky130_fd_sc_hd__or2_1 _5326_ (.A(net643),
    .B(net279),
    .X(_2719_));
 sky130_fd_sc_hd__o211a_1 _5327_ (.A1(net2041),
    .A2(net295),
    .B1(net165),
    .C1(_2719_),
    .X(_0388_));
 sky130_fd_sc_hd__or2_1 _5328_ (.A(net884),
    .B(net282),
    .X(_2720_));
 sky130_fd_sc_hd__o211a_1 _5329_ (.A1(net2036),
    .A2(net299),
    .B1(net167),
    .C1(_2720_),
    .X(_0389_));
 sky130_fd_sc_hd__or2_1 _5330_ (.A(net835),
    .B(net279),
    .X(_2721_));
 sky130_fd_sc_hd__o211a_1 _5331_ (.A1(net2089),
    .A2(net297),
    .B1(net166),
    .C1(_2721_),
    .X(_0390_));
 sky130_fd_sc_hd__or2_1 _5332_ (.A(net845),
    .B(net277),
    .X(_2722_));
 sky130_fd_sc_hd__o211a_1 _5333_ (.A1(net2077),
    .A2(net296),
    .B1(net166),
    .C1(_2722_),
    .X(_0391_));
 sky130_fd_sc_hd__or2_1 _5334_ (.A(net843),
    .B(net283),
    .X(_2723_));
 sky130_fd_sc_hd__o211a_1 _5335_ (.A1(net2081),
    .A2(net299),
    .B1(net167),
    .C1(_2723_),
    .X(_0392_));
 sky130_fd_sc_hd__or2_1 _5336_ (.A(net689),
    .B(net283),
    .X(_2724_));
 sky130_fd_sc_hd__o211a_1 _5337_ (.A1(net2071),
    .A2(net299),
    .B1(net167),
    .C1(_2724_),
    .X(_0393_));
 sky130_fd_sc_hd__or2_1 _5338_ (.A(net1034),
    .B(net285),
    .X(_2725_));
 sky130_fd_sc_hd__o211a_1 _5339_ (.A1(net2104),
    .A2(net300),
    .B1(net167),
    .C1(_2725_),
    .X(_0394_));
 sky130_fd_sc_hd__or2_1 _5340_ (.A(net625),
    .B(net285),
    .X(_2726_));
 sky130_fd_sc_hd__o211a_1 _5341_ (.A1(net2068),
    .A2(net300),
    .B1(net169),
    .C1(_2726_),
    .X(_0395_));
 sky130_fd_sc_hd__or2_1 _5342_ (.A(net701),
    .B(net283),
    .X(_2727_));
 sky130_fd_sc_hd__o211a_1 _5343_ (.A1(net2069),
    .A2(net299),
    .B1(net167),
    .C1(_2727_),
    .X(_0396_));
 sky130_fd_sc_hd__or2_1 _5344_ (.A(net1096),
    .B(net284),
    .X(_2728_));
 sky130_fd_sc_hd__o211a_1 _5345_ (.A1(net2096),
    .A2(net299),
    .B1(net167),
    .C1(_2728_),
    .X(_0397_));
 sky130_fd_sc_hd__or2_1 _5346_ (.A(net880),
    .B(net289),
    .X(_2729_));
 sky130_fd_sc_hd__o211a_1 _5347_ (.A1(net2051),
    .A2(net302),
    .B1(net168),
    .C1(_2729_),
    .X(_0398_));
 sky130_fd_sc_hd__or2_1 _5348_ (.A(net859),
    .B(net286),
    .X(_2730_));
 sky130_fd_sc_hd__o211a_1 _5349_ (.A1(net2116),
    .A2(net300),
    .B1(net169),
    .C1(_2730_),
    .X(_0399_));
 sky130_fd_sc_hd__or2_1 _5350_ (.A(net976),
    .B(net274),
    .X(_2731_));
 sky130_fd_sc_hd__o211a_1 _5351_ (.A1(net2080),
    .A2(net293),
    .B1(net164),
    .C1(_2731_),
    .X(_0400_));
 sky130_fd_sc_hd__or2_1 _5352_ (.A(net956),
    .B(net276),
    .X(_2732_));
 sky130_fd_sc_hd__o211a_1 _5353_ (.A1(net2090),
    .A2(net294),
    .B1(net164),
    .C1(_2732_),
    .X(_0401_));
 sky130_fd_sc_hd__or2_1 _5354_ (.A(net1026),
    .B(net287),
    .X(_2733_));
 sky130_fd_sc_hd__o211a_1 _5355_ (.A1(net2083),
    .A2(net303),
    .B1(net169),
    .C1(_2733_),
    .X(_0402_));
 sky130_fd_sc_hd__or2_1 _5356_ (.A(net912),
    .B(net274),
    .X(_2734_));
 sky130_fd_sc_hd__o211a_1 _5357_ (.A1(net2064),
    .A2(net293),
    .B1(net164),
    .C1(_2734_),
    .X(_0403_));
 sky130_fd_sc_hd__or2_1 _5358_ (.A(net1048),
    .B(net280),
    .X(_2735_));
 sky130_fd_sc_hd__o211a_1 _5359_ (.A1(net2088),
    .A2(net298),
    .B1(net170),
    .C1(_2735_),
    .X(_0404_));
 sky130_fd_sc_hd__or2_1 _5360_ (.A(net1140),
    .B(net274),
    .X(_2736_));
 sky130_fd_sc_hd__o211a_1 _5361_ (.A1(net2075),
    .A2(net293),
    .B1(net164),
    .C1(_2736_),
    .X(_0405_));
 sky130_fd_sc_hd__or2_1 _5362_ (.A(net1208),
    .B(net275),
    .X(_2737_));
 sky130_fd_sc_hd__o211a_1 _5363_ (.A1(net2102),
    .A2(net293),
    .B1(net164),
    .C1(_2737_),
    .X(_0406_));
 sky130_fd_sc_hd__or2_1 _5364_ (.A(net1210),
    .B(net281),
    .X(_2738_));
 sky130_fd_sc_hd__o211a_1 _5365_ (.A1(net2095),
    .A2(net294),
    .B1(net164),
    .C1(_2738_),
    .X(_0407_));
 sky130_fd_sc_hd__or2_1 _5366_ (.A(net926),
    .B(net272),
    .X(_2739_));
 sky130_fd_sc_hd__o211a_1 _5367_ (.A1(net2076),
    .A2(net295),
    .B1(net165),
    .C1(_2739_),
    .X(_0408_));
 sky130_fd_sc_hd__or2_1 _5368_ (.A(net817),
    .B(net272),
    .X(_2740_));
 sky130_fd_sc_hd__o211a_1 _5369_ (.A1(net2097),
    .A2(net295),
    .B1(net165),
    .C1(_2740_),
    .X(_0409_));
 sky130_fd_sc_hd__or2_1 _5370_ (.A(net1170),
    .B(net273),
    .X(_2741_));
 sky130_fd_sc_hd__o211a_1 _5371_ (.A1(net2082),
    .A2(net295),
    .B1(net165),
    .C1(_2741_),
    .X(_0410_));
 sky130_fd_sc_hd__or2_1 _5372_ (.A(net962),
    .B(net280),
    .X(_2742_));
 sky130_fd_sc_hd__o211a_1 _5373_ (.A1(net2078),
    .A2(net298),
    .B1(net170),
    .C1(_2742_),
    .X(_0411_));
 sky130_fd_sc_hd__or2_4 _5374_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .X(_2743_));
 sky130_fd_sc_hd__o311ai_4 _5375_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .A2(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .A3(_2743_),
    .B1(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .C1(net469),
    .Y(_2744_));
 sky130_fd_sc_hd__nand2_1 _5376_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .Y(_2745_));
 sky130_fd_sc_hd__nor2_1 _5377_ (.A(_2744_),
    .B(_2745_),
    .Y(_2746_));
 sky130_fd_sc_hd__or2_4 _5378_ (.A(_2744_),
    .B(_2745_),
    .X(_2747_));
 sky130_fd_sc_hd__and3_4 _5379_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(_1412_),
    .C(_2746_),
    .X(_2748_));
 sky130_fd_sc_hd__or3_2 _5380_ (.A(_1411_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .C(_2747_),
    .X(_2749_));
 sky130_fd_sc_hd__nor2_4 _5381_ (.A(net473),
    .B(net270),
    .Y(_2750_));
 sky130_fd_sc_hd__nand2_1 _5382_ (.A(net469),
    .B(_2749_),
    .Y(_2751_));
 sky130_fd_sc_hd__o22a_1 _5383_ (.A1(net331),
    .A2(_2749_),
    .B1(_2751_),
    .B2(net1695),
    .X(_0412_));
 sky130_fd_sc_hd__a22o_1 _5384_ (.A1(net332),
    .A2(net271),
    .B1(net237),
    .B2(net1194),
    .X(_0413_));
 sky130_fd_sc_hd__o22a_1 _5385_ (.A1(net333),
    .A2(_2749_),
    .B1(_2751_),
    .B2(net900),
    .X(_0414_));
 sky130_fd_sc_hd__o22a_1 _5386_ (.A1(net334),
    .A2(_2749_),
    .B1(_2751_),
    .B2(net892),
    .X(_0415_));
 sky130_fd_sc_hd__a22o_1 _5387_ (.A1(net329),
    .A2(net271),
    .B1(net237),
    .B2(net1154),
    .X(_0416_));
 sky130_fd_sc_hd__a22o_1 _5388_ (.A1(_1741_),
    .A2(net271),
    .B1(net237),
    .B2(net1148),
    .X(_0417_));
 sky130_fd_sc_hd__a22o_1 _5389_ (.A1(net328),
    .A2(net271),
    .B1(net237),
    .B2(net1724),
    .X(_0418_));
 sky130_fd_sc_hd__a22o_1 _5390_ (.A1(net330),
    .A2(net270),
    .B1(net236),
    .B2(net1062),
    .X(_0419_));
 sky130_fd_sc_hd__a22o_1 _5391_ (.A1(net325),
    .A2(net270),
    .B1(net236),
    .B2(net1270),
    .X(_0420_));
 sky130_fd_sc_hd__a22o_1 _5392_ (.A1(net327),
    .A2(net271),
    .B1(net237),
    .B2(net1030),
    .X(_0421_));
 sky130_fd_sc_hd__a22o_1 _5393_ (.A1(net326),
    .A2(net270),
    .B1(net236),
    .B2(net1559),
    .X(_0422_));
 sky130_fd_sc_hd__a22o_1 _5394_ (.A1(net324),
    .A2(net270),
    .B1(net236),
    .B2(net1623),
    .X(_0423_));
 sky130_fd_sc_hd__a22o_1 _5395_ (.A1(net321),
    .A2(net271),
    .B1(net237),
    .B2(net1142),
    .X(_0424_));
 sky130_fd_sc_hd__a22o_1 _5396_ (.A1(net323),
    .A2(net271),
    .B1(net237),
    .B2(net1573),
    .X(_0425_));
 sky130_fd_sc_hd__a22o_1 _5397_ (.A1(net322),
    .A2(net271),
    .B1(net237),
    .B2(net1457),
    .X(_0426_));
 sky130_fd_sc_hd__a22o_1 _5398_ (.A1(net320),
    .A2(net271),
    .B1(net237),
    .B2(net1599),
    .X(_0427_));
 sky130_fd_sc_hd__a22o_1 _5399_ (.A1(net344),
    .A2(net270),
    .B1(net236),
    .B2(net1070),
    .X(_0428_));
 sky130_fd_sc_hd__a22o_1 _5400_ (.A1(_1512_),
    .A2(net271),
    .B1(net236),
    .B2(net1712),
    .X(_0429_));
 sky130_fd_sc_hd__a22o_1 _5401_ (.A1(net343),
    .A2(net271),
    .B1(net237),
    .B2(net1503),
    .X(_0430_));
 sky130_fd_sc_hd__a22o_1 _5402_ (.A1(net345),
    .A2(net271),
    .B1(net237),
    .B2(net1032),
    .X(_0431_));
 sky130_fd_sc_hd__a22o_1 _5403_ (.A1(net340),
    .A2(net270),
    .B1(net236),
    .B2(net1084),
    .X(_0432_));
 sky130_fd_sc_hd__a22o_1 _5404_ (.A1(net342),
    .A2(net270),
    .B1(net236),
    .B2(net968),
    .X(_0433_));
 sky130_fd_sc_hd__a22o_1 _5405_ (.A1(net341),
    .A2(net271),
    .B1(net237),
    .B2(net1693),
    .X(_0434_));
 sky130_fd_sc_hd__a22o_1 _5406_ (.A1(net339),
    .A2(net270),
    .B1(net236),
    .B2(net1641),
    .X(_0435_));
 sky130_fd_sc_hd__a22o_1 _5407_ (.A1(net336),
    .A2(net271),
    .B1(net237),
    .B2(net1509),
    .X(_0436_));
 sky130_fd_sc_hd__a22o_1 _5408_ (.A1(net338),
    .A2(net270),
    .B1(net236),
    .B2(net1603),
    .X(_0437_));
 sky130_fd_sc_hd__a22o_1 _5409_ (.A1(net337),
    .A2(net270),
    .B1(net236),
    .B2(net1186),
    .X(_0438_));
 sky130_fd_sc_hd__a22o_1 _5410_ (.A1(net335),
    .A2(net270),
    .B1(net236),
    .B2(net1527),
    .X(_0439_));
 sky130_fd_sc_hd__a22o_1 _5411_ (.A1(net348),
    .A2(net270),
    .B1(net236),
    .B2(net1625),
    .X(_0440_));
 sky130_fd_sc_hd__a22o_1 _5412_ (.A1(net346),
    .A2(net270),
    .B1(net236),
    .B2(net1102),
    .X(_0441_));
 sky130_fd_sc_hd__a22o_1 _5413_ (.A1(net347),
    .A2(net270),
    .B1(net236),
    .B2(net1325),
    .X(_0442_));
 sky130_fd_sc_hd__a22o_1 _5414_ (.A1(net370),
    .A2(net270),
    .B1(net236),
    .B2(net1040),
    .X(_0443_));
 sky130_fd_sc_hd__or3_4 _5415_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(_1412_),
    .C(_2744_),
    .X(_2752_));
 sky130_fd_sc_hd__nand2_2 _5416_ (.A(_1413_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .Y(_2753_));
 sky130_fd_sc_hd__nor2_4 _5417_ (.A(_2752_),
    .B(_2753_),
    .Y(_2754_));
 sky130_fd_sc_hd__or2_1 _5418_ (.A(_2752_),
    .B(_2753_),
    .X(_2755_));
 sky130_fd_sc_hd__nor2_4 _5419_ (.A(net473),
    .B(net268),
    .Y(_2756_));
 sky130_fd_sc_hd__nand2_1 _5420_ (.A(net467),
    .B(_2755_),
    .Y(_2757_));
 sky130_fd_sc_hd__a22o_1 _5421_ (.A1(net331),
    .A2(net269),
    .B1(net235),
    .B2(net990),
    .X(_0444_));
 sky130_fd_sc_hd__o22a_1 _5422_ (.A1(net332),
    .A2(_2755_),
    .B1(_2757_),
    .B2(net908),
    .X(_0445_));
 sky130_fd_sc_hd__a22o_1 _5423_ (.A1(net333),
    .A2(net269),
    .B1(net235),
    .B2(net1673),
    .X(_0446_));
 sky130_fd_sc_hd__o22a_1 _5424_ (.A1(net334),
    .A2(_2755_),
    .B1(_2757_),
    .B2(net1138),
    .X(_0447_));
 sky130_fd_sc_hd__a22o_1 _5425_ (.A1(net329),
    .A2(net269),
    .B1(net235),
    .B2(net1246),
    .X(_0448_));
 sky130_fd_sc_hd__a22o_1 _5426_ (.A1(_1741_),
    .A2(net269),
    .B1(net235),
    .B2(net1150),
    .X(_0449_));
 sky130_fd_sc_hd__a22o_1 _5427_ (.A1(net328),
    .A2(net269),
    .B1(net234),
    .B2(net1611),
    .X(_0450_));
 sky130_fd_sc_hd__a22o_1 _5428_ (.A1(net330),
    .A2(net268),
    .B1(net234),
    .B2(net1451),
    .X(_0451_));
 sky130_fd_sc_hd__a22o_1 _5429_ (.A1(net325),
    .A2(net268),
    .B1(net234),
    .B2(net1074),
    .X(_0452_));
 sky130_fd_sc_hd__a22o_1 _5430_ (.A1(net327),
    .A2(net269),
    .B1(net235),
    .B2(net1252),
    .X(_0453_));
 sky130_fd_sc_hd__a22o_1 _5431_ (.A1(net326),
    .A2(net268),
    .B1(net234),
    .B2(net1244),
    .X(_0454_));
 sky130_fd_sc_hd__a22o_1 _5432_ (.A1(net324),
    .A2(net268),
    .B1(net234),
    .B2(net1262),
    .X(_0455_));
 sky130_fd_sc_hd__a22o_1 _5433_ (.A1(net321),
    .A2(net269),
    .B1(net235),
    .B2(net1401),
    .X(_0456_));
 sky130_fd_sc_hd__a22o_1 _5434_ (.A1(net323),
    .A2(net269),
    .B1(net235),
    .B2(net1216),
    .X(_0457_));
 sky130_fd_sc_hd__a22o_1 _5435_ (.A1(net322),
    .A2(net269),
    .B1(net235),
    .B2(net1541),
    .X(_0458_));
 sky130_fd_sc_hd__a22o_1 _5436_ (.A1(net320),
    .A2(net269),
    .B1(net235),
    .B2(net1168),
    .X(_0459_));
 sky130_fd_sc_hd__a22o_1 _5437_ (.A1(net344),
    .A2(net268),
    .B1(net234),
    .B2(net1220),
    .X(_0460_));
 sky130_fd_sc_hd__a22o_1 _5438_ (.A1(_1512_),
    .A2(net269),
    .B1(net235),
    .B2(net1353),
    .X(_0461_));
 sky130_fd_sc_hd__a22o_1 _5439_ (.A1(net343),
    .A2(net269),
    .B1(net235),
    .B2(net1104),
    .X(_0462_));
 sky130_fd_sc_hd__a22o_1 _5440_ (.A1(net345),
    .A2(net269),
    .B1(net235),
    .B2(net1110),
    .X(_0463_));
 sky130_fd_sc_hd__a22o_1 _5441_ (.A1(net340),
    .A2(net268),
    .B1(net234),
    .B2(net996),
    .X(_0464_));
 sky130_fd_sc_hd__a22o_1 _5442_ (.A1(net342),
    .A2(net268),
    .B1(net234),
    .B2(net1024),
    .X(_0465_));
 sky130_fd_sc_hd__a22o_1 _5443_ (.A1(net341),
    .A2(net269),
    .B1(net235),
    .B2(net1184),
    .X(_0466_));
 sky130_fd_sc_hd__a22o_1 _5444_ (.A1(net339),
    .A2(net268),
    .B1(net234),
    .B2(net1551),
    .X(_0467_));
 sky130_fd_sc_hd__a22o_1 _5445_ (.A1(net336),
    .A2(net269),
    .B1(net235),
    .B2(net1046),
    .X(_0468_));
 sky130_fd_sc_hd__a22o_1 _5446_ (.A1(net338),
    .A2(net268),
    .B1(net234),
    .B2(net1301),
    .X(_0469_));
 sky130_fd_sc_hd__a22o_1 _5447_ (.A1(net337),
    .A2(net268),
    .B1(net234),
    .B2(net984),
    .X(_0470_));
 sky130_fd_sc_hd__a22o_1 _5448_ (.A1(net335),
    .A2(net268),
    .B1(net234),
    .B2(net1258),
    .X(_0471_));
 sky130_fd_sc_hd__a22o_1 _5449_ (.A1(net348),
    .A2(net268),
    .B1(net234),
    .B2(net1403),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _5450_ (.A1(net346),
    .A2(net268),
    .B1(net234),
    .B2(net1042),
    .X(_0473_));
 sky130_fd_sc_hd__a22o_1 _5451_ (.A1(net347),
    .A2(net268),
    .B1(net234),
    .B2(net1431),
    .X(_0474_));
 sky130_fd_sc_hd__a22o_1 _5452_ (.A1(net370),
    .A2(net268),
    .B1(net234),
    .B2(net1645),
    .X(_0475_));
 sky130_fd_sc_hd__or3_4 _5453_ (.A(_1411_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .C(net365),
    .X(_2758_));
 sky130_fd_sc_hd__nor2_1 _5454_ (.A(_2753_),
    .B(_2758_),
    .Y(_2759_));
 sky130_fd_sc_hd__or2_1 _5455_ (.A(_2753_),
    .B(_2758_),
    .X(_2760_));
 sky130_fd_sc_hd__nor2_1 _5456_ (.A(net479),
    .B(net266),
    .Y(_2761_));
 sky130_fd_sc_hd__nand2_1 _5457_ (.A(net467),
    .B(_2760_),
    .Y(_2762_));
 sky130_fd_sc_hd__o22a_1 _5458_ (.A1(net331),
    .A2(_2760_),
    .B1(_2762_),
    .B2(net855),
    .X(_0476_));
 sky130_fd_sc_hd__a22o_1 _5459_ (.A1(net332),
    .A2(net266),
    .B1(net233),
    .B2(net1280),
    .X(_0477_));
 sky130_fd_sc_hd__a22o_1 _5460_ (.A1(net333),
    .A2(net266),
    .B1(net233),
    .B2(net1393),
    .X(_0478_));
 sky130_fd_sc_hd__o22a_1 _5461_ (.A1(net334),
    .A2(_2760_),
    .B1(_2762_),
    .B2(net861),
    .X(_0479_));
 sky130_fd_sc_hd__a22o_1 _5462_ (.A1(net329),
    .A2(net266),
    .B1(net233),
    .B2(net1329),
    .X(_0480_));
 sky130_fd_sc_hd__a22o_1 _5463_ (.A1(_1741_),
    .A2(net266),
    .B1(net233),
    .B2(net1565),
    .X(_0481_));
 sky130_fd_sc_hd__a22o_1 _5464_ (.A1(net328),
    .A2(net266),
    .B1(net232),
    .B2(net1697),
    .X(_0482_));
 sky130_fd_sc_hd__a22o_1 _5465_ (.A1(net330),
    .A2(net267),
    .B1(net232),
    .B2(net1090),
    .X(_0483_));
 sky130_fd_sc_hd__a22o_1 _5466_ (.A1(net325),
    .A2(net267),
    .B1(net232),
    .B2(net948),
    .X(_0484_));
 sky130_fd_sc_hd__a22o_1 _5467_ (.A1(net327),
    .A2(net267),
    .B1(net233),
    .B2(net1513),
    .X(_0485_));
 sky130_fd_sc_hd__a22o_1 _5468_ (.A1(net326),
    .A2(net267),
    .B1(net232),
    .B2(net1601),
    .X(_0486_));
 sky130_fd_sc_hd__a22o_1 _5469_ (.A1(net324),
    .A2(net267),
    .B1(net232),
    .B2(net934),
    .X(_0487_));
 sky130_fd_sc_hd__a22o_1 _5470_ (.A1(net321),
    .A2(net266),
    .B1(net233),
    .B2(net1736),
    .X(_0488_));
 sky130_fd_sc_hd__a22o_1 _5471_ (.A1(net323),
    .A2(net266),
    .B1(net233),
    .B2(net1313),
    .X(_0489_));
 sky130_fd_sc_hd__a22o_1 _5472_ (.A1(net322),
    .A2(net266),
    .B1(net233),
    .B2(net1575),
    .X(_0490_));
 sky130_fd_sc_hd__a22o_1 _5473_ (.A1(net320),
    .A2(net266),
    .B1(net233),
    .B2(net1124),
    .X(_0491_));
 sky130_fd_sc_hd__a22o_1 _5474_ (.A1(net344),
    .A2(net267),
    .B1(net232),
    .B2(net1501),
    .X(_0492_));
 sky130_fd_sc_hd__a22o_1 _5475_ (.A1(_1512_),
    .A2(net266),
    .B1(net233),
    .B2(net1756),
    .X(_0493_));
 sky130_fd_sc_hd__a22o_1 _5476_ (.A1(net343),
    .A2(net266),
    .B1(net233),
    .B2(net1663),
    .X(_0494_));
 sky130_fd_sc_hd__a22o_1 _5477_ (.A1(net345),
    .A2(net266),
    .B1(net233),
    .B2(net1202),
    .X(_0495_));
 sky130_fd_sc_hd__a22o_1 _5478_ (.A1(net340),
    .A2(net267),
    .B1(net232),
    .B2(net1248),
    .X(_0496_));
 sky130_fd_sc_hd__a22o_1 _5479_ (.A1(net342),
    .A2(net267),
    .B1(net232),
    .B2(net1176),
    .X(_0497_));
 sky130_fd_sc_hd__a22o_1 _5480_ (.A1(net341),
    .A2(net266),
    .B1(net233),
    .B2(net1441),
    .X(_0498_));
 sky130_fd_sc_hd__a22o_1 _5481_ (.A1(net339),
    .A2(net267),
    .B1(net232),
    .B2(net1188),
    .X(_0499_));
 sky130_fd_sc_hd__a22o_1 _5482_ (.A1(net336),
    .A2(net266),
    .B1(net233),
    .B2(net1726),
    .X(_0500_));
 sky130_fd_sc_hd__a22o_1 _5483_ (.A1(net338),
    .A2(net267),
    .B1(net232),
    .B2(net1415),
    .X(_0501_));
 sky130_fd_sc_hd__a22o_1 _5484_ (.A1(net337),
    .A2(net267),
    .B1(net232),
    .B2(net1078),
    .X(_0502_));
 sky130_fd_sc_hd__a22o_1 _5485_ (.A1(net335),
    .A2(net266),
    .B1(net232),
    .B2(net1288),
    .X(_0503_));
 sky130_fd_sc_hd__a22o_1 _5486_ (.A1(net348),
    .A2(net267),
    .B1(net232),
    .B2(net1260),
    .X(_0504_));
 sky130_fd_sc_hd__a22o_1 _5487_ (.A1(net346),
    .A2(net267),
    .B1(net232),
    .B2(net1361),
    .X(_0505_));
 sky130_fd_sc_hd__a22o_1 _5488_ (.A1(net347),
    .A2(net267),
    .B1(net232),
    .B2(net1619),
    .X(_0506_));
 sky130_fd_sc_hd__a22o_1 _5489_ (.A1(net370),
    .A2(net267),
    .B1(net232),
    .B2(net1305),
    .X(_0507_));
 sky130_fd_sc_hd__and3_4 _5490_ (.A(_1411_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .C(_2746_),
    .X(_2763_));
 sky130_fd_sc_hd__or3_2 _5491_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(_1412_),
    .C(_2747_),
    .X(_2764_));
 sky130_fd_sc_hd__nor2_4 _5492_ (.A(net473),
    .B(net264),
    .Y(_2765_));
 sky130_fd_sc_hd__nand2_1 _5493_ (.A(net469),
    .B(_2764_),
    .Y(_2766_));
 sky130_fd_sc_hd__a22o_1 _5494_ (.A1(net331),
    .A2(net265),
    .B1(net231),
    .B2(net1264),
    .X(_0508_));
 sky130_fd_sc_hd__o22a_1 _5495_ (.A1(net332),
    .A2(_2764_),
    .B1(_2766_),
    .B2(net904),
    .X(_0509_));
 sky130_fd_sc_hd__o22a_1 _5496_ (.A1(net333),
    .A2(_2764_),
    .B1(_2766_),
    .B2(net982),
    .X(_0510_));
 sky130_fd_sc_hd__o22a_1 _5497_ (.A1(net334),
    .A2(_2764_),
    .B1(_2766_),
    .B2(net970),
    .X(_0511_));
 sky130_fd_sc_hd__a22o_1 _5498_ (.A1(net329),
    .A2(net265),
    .B1(net231),
    .B2(net1433),
    .X(_0512_));
 sky130_fd_sc_hd__a22o_1 _5499_ (.A1(_1741_),
    .A2(net265),
    .B1(net231),
    .B2(net1236),
    .X(_0513_));
 sky130_fd_sc_hd__a22o_1 _5500_ (.A1(net328),
    .A2(net265),
    .B1(net231),
    .B2(net1653),
    .X(_0514_));
 sky130_fd_sc_hd__a22o_1 _5501_ (.A1(net330),
    .A2(net264),
    .B1(net230),
    .B2(net1563),
    .X(_0515_));
 sky130_fd_sc_hd__a22o_1 _5502_ (.A1(net325),
    .A2(net264),
    .B1(net230),
    .B2(net1497),
    .X(_0516_));
 sky130_fd_sc_hd__a22o_1 _5503_ (.A1(net327),
    .A2(net265),
    .B1(net231),
    .B2(net1144),
    .X(_0517_));
 sky130_fd_sc_hd__a22o_1 _5504_ (.A1(net326),
    .A2(net264),
    .B1(net230),
    .B2(net1254),
    .X(_0518_));
 sky130_fd_sc_hd__a22o_1 _5505_ (.A1(net324),
    .A2(net264),
    .B1(net230),
    .B2(net1561),
    .X(_0519_));
 sky130_fd_sc_hd__a22o_1 _5506_ (.A1(net321),
    .A2(net265),
    .B1(net231),
    .B2(net940),
    .X(_0520_));
 sky130_fd_sc_hd__a22o_1 _5507_ (.A1(net323),
    .A2(net265),
    .B1(net231),
    .B2(net1591),
    .X(_0521_));
 sky130_fd_sc_hd__a22o_1 _5508_ (.A1(net322),
    .A2(net265),
    .B1(net231),
    .B2(net1349),
    .X(_0522_));
 sky130_fd_sc_hd__a22o_1 _5509_ (.A1(net320),
    .A2(net265),
    .B1(net231),
    .B2(net1190),
    .X(_0523_));
 sky130_fd_sc_hd__a22o_1 _5510_ (.A1(net344),
    .A2(net264),
    .B1(net230),
    .B2(net1447),
    .X(_0524_));
 sky130_fd_sc_hd__a22o_1 _5511_ (.A1(_1512_),
    .A2(net265),
    .B1(net230),
    .B2(net1555),
    .X(_0525_));
 sky130_fd_sc_hd__a22o_1 _5512_ (.A1(net343),
    .A2(net265),
    .B1(net231),
    .B2(net1036),
    .X(_0526_));
 sky130_fd_sc_hd__a22o_1 _5513_ (.A1(net345),
    .A2(net265),
    .B1(net231),
    .B2(net1477),
    .X(_0527_));
 sky130_fd_sc_hd__a22o_1 _5514_ (.A1(net340),
    .A2(net264),
    .B1(net230),
    .B2(net1303),
    .X(_0528_));
 sky130_fd_sc_hd__a22o_1 _5515_ (.A1(net342),
    .A2(net264),
    .B1(net230),
    .B2(net1008),
    .X(_0529_));
 sky130_fd_sc_hd__a22o_1 _5516_ (.A1(net341),
    .A2(net265),
    .B1(net231),
    .B2(net1198),
    .X(_0530_));
 sky130_fd_sc_hd__a22o_1 _5517_ (.A1(net339),
    .A2(net264),
    .B1(net230),
    .B2(net1537),
    .X(_0531_));
 sky130_fd_sc_hd__a22o_1 _5518_ (.A1(net336),
    .A2(net265),
    .B1(net231),
    .B2(net1397),
    .X(_0532_));
 sky130_fd_sc_hd__a22o_1 _5519_ (.A1(net338),
    .A2(net264),
    .B1(net230),
    .B2(net1064),
    .X(_0533_));
 sky130_fd_sc_hd__a22o_1 _5520_ (.A1(net337),
    .A2(net264),
    .B1(net230),
    .B2(net1082),
    .X(_0534_));
 sky130_fd_sc_hd__a22o_1 _5521_ (.A1(net335),
    .A2(net264),
    .B1(net230),
    .B2(net1579),
    .X(_0535_));
 sky130_fd_sc_hd__a22o_1 _5522_ (.A1(net348),
    .A2(net264),
    .B1(net230),
    .B2(net1250),
    .X(_0536_));
 sky130_fd_sc_hd__a22o_1 _5523_ (.A1(net346),
    .A2(net264),
    .B1(net230),
    .B2(net1439),
    .X(_0537_));
 sky130_fd_sc_hd__a22o_1 _5524_ (.A1(net347),
    .A2(net264),
    .B1(net230),
    .B2(net1615),
    .X(_0538_));
 sky130_fd_sc_hd__a22o_1 _5525_ (.A1(net370),
    .A2(net264),
    .B1(net230),
    .B2(net1238),
    .X(_0539_));
 sky130_fd_sc_hd__nand2_8 _5526_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .Y(_2767_));
 sky130_fd_sc_hd__nor2_8 _5527_ (.A(_2747_),
    .B(_2767_),
    .Y(_2768_));
 sky130_fd_sc_hd__or2_2 _5528_ (.A(_2747_),
    .B(_2767_),
    .X(_2769_));
 sky130_fd_sc_hd__nor2_4 _5529_ (.A(net473),
    .B(net262),
    .Y(_2770_));
 sky130_fd_sc_hd__nand2_2 _5530_ (.A(net469),
    .B(_2769_),
    .Y(_2771_));
 sky130_fd_sc_hd__o22a_1 _5531_ (.A1(net331),
    .A2(_2769_),
    .B1(_2771_),
    .B2(net1842),
    .X(_0540_));
 sky130_fd_sc_hd__o22a_1 _5532_ (.A1(net332),
    .A2(_2769_),
    .B1(_2771_),
    .B2(net866),
    .X(_0541_));
 sky130_fd_sc_hd__o22a_1 _5533_ (.A1(net333),
    .A2(_2769_),
    .B1(_2771_),
    .B2(net914),
    .X(_0542_));
 sky130_fd_sc_hd__o22a_1 _5534_ (.A1(net334),
    .A2(_2769_),
    .B1(_2771_),
    .B2(net872),
    .X(_0543_));
 sky130_fd_sc_hd__a22o_1 _5535_ (.A1(net329),
    .A2(net263),
    .B1(net229),
    .B2(net1228),
    .X(_0544_));
 sky130_fd_sc_hd__a22o_1 _5536_ (.A1(_1741_),
    .A2(net263),
    .B1(net229),
    .B2(net930),
    .X(_0545_));
 sky130_fd_sc_hd__a22o_1 _5537_ (.A1(net328),
    .A2(net263),
    .B1(net229),
    .B2(net1359),
    .X(_0546_));
 sky130_fd_sc_hd__a22o_1 _5538_ (.A1(net330),
    .A2(net262),
    .B1(net228),
    .B2(net1060),
    .X(_0547_));
 sky130_fd_sc_hd__a22o_1 _5539_ (.A1(net325),
    .A2(net262),
    .B1(net228),
    .B2(net1206),
    .X(_0548_));
 sky130_fd_sc_hd__a22o_1 _5540_ (.A1(net327),
    .A2(net263),
    .B1(net229),
    .B2(net1166),
    .X(_0549_));
 sky130_fd_sc_hd__a22o_1 _5541_ (.A1(net326),
    .A2(net262),
    .B1(net228),
    .B2(net1182),
    .X(_0550_));
 sky130_fd_sc_hd__a22o_1 _5542_ (.A1(net324),
    .A2(net262),
    .B1(net228),
    .B2(net1455),
    .X(_0551_));
 sky130_fd_sc_hd__a22o_1 _5543_ (.A1(net321),
    .A2(net263),
    .B1(net229),
    .B2(net1000),
    .X(_0552_));
 sky130_fd_sc_hd__a22o_1 _5544_ (.A1(net323),
    .A2(net263),
    .B1(net229),
    .B2(net1489),
    .X(_0553_));
 sky130_fd_sc_hd__a22o_1 _5545_ (.A1(net322),
    .A2(net263),
    .B1(net229),
    .B2(net1242),
    .X(_0554_));
 sky130_fd_sc_hd__a22o_1 _5546_ (.A1(net320),
    .A2(net263),
    .B1(net229),
    .B2(net1804),
    .X(_0555_));
 sky130_fd_sc_hd__a22o_1 _5547_ (.A1(net344),
    .A2(net262),
    .B1(net228),
    .B2(net1732),
    .X(_0556_));
 sky130_fd_sc_hd__a22o_1 _5548_ (.A1(_1512_),
    .A2(net263),
    .B1(net228),
    .B2(net1174),
    .X(_0557_));
 sky130_fd_sc_hd__a22o_1 _5549_ (.A1(net343),
    .A2(net263),
    .B1(net229),
    .B2(net1337),
    .X(_0558_));
 sky130_fd_sc_hd__a22o_1 _5550_ (.A1(net345),
    .A2(net263),
    .B1(net229),
    .B2(net1319),
    .X(_0559_));
 sky130_fd_sc_hd__a22o_1 _5551_ (.A1(net340),
    .A2(net262),
    .B1(net228),
    .B2(net1687),
    .X(_0560_));
 sky130_fd_sc_hd__a22o_1 _5552_ (.A1(net342),
    .A2(net262),
    .B1(net228),
    .B2(net1309),
    .X(_0561_));
 sky130_fd_sc_hd__a22o_1 _5553_ (.A1(net341),
    .A2(net263),
    .B1(net229),
    .B2(net1744),
    .X(_0562_));
 sky130_fd_sc_hd__a22o_1 _5554_ (.A1(net339),
    .A2(net262),
    .B1(net228),
    .B2(net1818),
    .X(_0563_));
 sky130_fd_sc_hd__a22o_1 _5555_ (.A1(net336),
    .A2(net263),
    .B1(net229),
    .B2(net1094),
    .X(_0564_));
 sky130_fd_sc_hd__a22o_1 _5556_ (.A1(net338),
    .A2(net262),
    .B1(net228),
    .B2(net1297),
    .X(_0565_));
 sky130_fd_sc_hd__a22o_1 _5557_ (.A1(net337),
    .A2(net262),
    .B1(net228),
    .B2(net1230),
    .X(_0566_));
 sky130_fd_sc_hd__a22o_1 _5558_ (.A1(net335),
    .A2(net262),
    .B1(net228),
    .B2(net1389),
    .X(_0567_));
 sky130_fd_sc_hd__a22o_1 _5559_ (.A1(net348),
    .A2(net262),
    .B1(net228),
    .B2(net1369),
    .X(_0568_));
 sky130_fd_sc_hd__a22o_1 _5560_ (.A1(net346),
    .A2(net262),
    .B1(net228),
    .B2(net988),
    .X(_0569_));
 sky130_fd_sc_hd__a22o_1 _5561_ (.A1(net347),
    .A2(net262),
    .B1(net228),
    .B2(net1453),
    .X(_0570_));
 sky130_fd_sc_hd__a22o_1 _5562_ (.A1(net370),
    .A2(net262),
    .B1(net228),
    .B2(net1519),
    .X(_0571_));
 sky130_fd_sc_hd__nor2_4 _5563_ (.A(_2743_),
    .B(_2747_),
    .Y(_2772_));
 sky130_fd_sc_hd__inv_2 _5564_ (.A(net260),
    .Y(_2773_));
 sky130_fd_sc_hd__nor2_4 _5565_ (.A(net479),
    .B(net260),
    .Y(_2774_));
 sky130_fd_sc_hd__or2_1 _5566_ (.A(net480),
    .B(net260),
    .X(_2775_));
 sky130_fd_sc_hd__a22o_1 _5567_ (.A1(net331),
    .A2(net260),
    .B1(net227),
    .B2(net1180),
    .X(_0572_));
 sky130_fd_sc_hd__a22o_1 _5568_ (.A1(net332),
    .A2(net260),
    .B1(net227),
    .B2(net1720),
    .X(_0573_));
 sky130_fd_sc_hd__o22a_1 _5569_ (.A1(net333),
    .A2(_2773_),
    .B1(_2775_),
    .B2(net1022),
    .X(_0574_));
 sky130_fd_sc_hd__o22a_1 _5570_ (.A1(net334),
    .A2(_2773_),
    .B1(_2775_),
    .B2(net1413),
    .X(_0575_));
 sky130_fd_sc_hd__a22o_1 _5571_ (.A1(net329),
    .A2(net260),
    .B1(net227),
    .B2(net1679),
    .X(_0576_));
 sky130_fd_sc_hd__a22o_1 _5572_ (.A1(_1741_),
    .A2(net260),
    .B1(net227),
    .B2(net1683),
    .X(_0577_));
 sky130_fd_sc_hd__a22o_1 _5573_ (.A1(net328),
    .A2(net260),
    .B1(net226),
    .B2(net1677),
    .X(_0578_));
 sky130_fd_sc_hd__a22o_1 _5574_ (.A1(net330),
    .A2(net261),
    .B1(net226),
    .B2(net1429),
    .X(_0579_));
 sky130_fd_sc_hd__a22o_1 _5575_ (.A1(net325),
    .A2(net261),
    .B1(net226),
    .B2(net1367),
    .X(_0580_));
 sky130_fd_sc_hd__a22o_1 _5576_ (.A1(net327),
    .A2(net260),
    .B1(net227),
    .B2(net1547),
    .X(_0581_));
 sky130_fd_sc_hd__a22o_1 _5577_ (.A1(net326),
    .A2(net261),
    .B1(net226),
    .B2(net1479),
    .X(_0582_));
 sky130_fd_sc_hd__a22o_1 _5578_ (.A1(net324),
    .A2(net261),
    .B1(net226),
    .B2(net1387),
    .X(_0583_));
 sky130_fd_sc_hd__a22o_1 _5579_ (.A1(net321),
    .A2(net260),
    .B1(net227),
    .B2(net1391),
    .X(_0584_));
 sky130_fd_sc_hd__a22o_1 _5580_ (.A1(net323),
    .A2(_2772_),
    .B1(net227),
    .B2(net1553),
    .X(_0585_));
 sky130_fd_sc_hd__a22o_1 _5581_ (.A1(net322),
    .A2(_2772_),
    .B1(net227),
    .B2(net1437),
    .X(_0586_));
 sky130_fd_sc_hd__a22o_1 _5582_ (.A1(net320),
    .A2(net260),
    .B1(net227),
    .B2(net1493),
    .X(_0587_));
 sky130_fd_sc_hd__a22o_1 _5583_ (.A1(net344),
    .A2(net261),
    .B1(net226),
    .B2(net1703),
    .X(_0588_));
 sky130_fd_sc_hd__a22o_1 _5584_ (.A1(_1512_),
    .A2(net260),
    .B1(net227),
    .B2(net1794),
    .X(_0589_));
 sky130_fd_sc_hd__a22o_1 _5585_ (.A1(net343),
    .A2(net260),
    .B1(net227),
    .B2(net986),
    .X(_0590_));
 sky130_fd_sc_hd__a22o_1 _5586_ (.A1(net345),
    .A2(net260),
    .B1(net227),
    .B2(net1214),
    .X(_0591_));
 sky130_fd_sc_hd__a22o_1 _5587_ (.A1(_1584_),
    .A2(net261),
    .B1(net226),
    .B2(net1587),
    .X(_0592_));
 sky130_fd_sc_hd__a22o_1 _5588_ (.A1(net342),
    .A2(net261),
    .B1(net226),
    .B2(net1056),
    .X(_0593_));
 sky130_fd_sc_hd__a22o_1 _5589_ (.A1(net341),
    .A2(net260),
    .B1(net227),
    .B2(net1491),
    .X(_0594_));
 sky130_fd_sc_hd__a22o_1 _5590_ (.A1(net339),
    .A2(net261),
    .B1(net226),
    .B2(net1824),
    .X(_0595_));
 sky130_fd_sc_hd__a22o_1 _5591_ (.A1(net336),
    .A2(net260),
    .B1(net227),
    .B2(net1647),
    .X(_0596_));
 sky130_fd_sc_hd__a22o_1 _5592_ (.A1(_1607_),
    .A2(net261),
    .B1(net226),
    .B2(net1740),
    .X(_0597_));
 sky130_fd_sc_hd__a22o_1 _5593_ (.A1(net337),
    .A2(net261),
    .B1(net226),
    .B2(net1224),
    .X(_0598_));
 sky130_fd_sc_hd__a22o_1 _5594_ (.A1(net335),
    .A2(net261),
    .B1(net226),
    .B2(net1657),
    .X(_0599_));
 sky130_fd_sc_hd__a22o_1 _5595_ (.A1(net348),
    .A2(net261),
    .B1(net226),
    .B2(net1691),
    .X(_0600_));
 sky130_fd_sc_hd__a22o_1 _5596_ (.A1(net346),
    .A2(net261),
    .B1(net226),
    .B2(net1681),
    .X(_0601_));
 sky130_fd_sc_hd__a22o_1 _5597_ (.A1(net347),
    .A2(net261),
    .B1(net226),
    .B2(net1395),
    .X(_0602_));
 sky130_fd_sc_hd__a22o_1 _5598_ (.A1(net370),
    .A2(net261),
    .B1(net226),
    .B2(net1649),
    .X(_0603_));
 sky130_fd_sc_hd__and2_4 _5599_ (.A(net175),
    .B(net279),
    .X(_2776_));
 sky130_fd_sc_hd__nand2_1 _5600_ (.A(net179),
    .B(net284),
    .Y(_2777_));
 sky130_fd_sc_hd__o31ai_1 _5601_ (.A1(net2194),
    .A2(net2203),
    .A3(_2267_),
    .B1(net2059),
    .Y(_2778_));
 sky130_fd_sc_hd__or3b_1 _5602_ (.A(_2267_),
    .B(net2194),
    .C_N(net2203),
    .X(_2779_));
 sky130_fd_sc_hd__nor2_1 _5603_ (.A(net2197),
    .B(_2779_),
    .Y(_2780_));
 sky130_fd_sc_hd__nor2_1 _5604_ (.A(net2058),
    .B(_2263_),
    .Y(_2781_));
 sky130_fd_sc_hd__nor2_1 _5605_ (.A(net2197),
    .B(net2203),
    .Y(_2782_));
 sky130_fd_sc_hd__a41o_1 _5606_ (.A1(_1407_),
    .A2(net2058),
    .A3(net2073),
    .A4(_2782_),
    .B1(_2780_),
    .X(_2783_));
 sky130_fd_sc_hd__o31a_1 _5607_ (.A1(_2778_),
    .A2(_2781_),
    .A3(_2783_),
    .B1(_2776_),
    .X(_0604_));
 sky130_fd_sc_hd__nor3_1 _5608_ (.A(net2055),
    .B(net2092),
    .C(net2010),
    .Y(_2784_));
 sky130_fd_sc_hd__a21oi_2 _5609_ (.A1(net2197),
    .A2(_2784_),
    .B1(_2779_),
    .Y(_2785_));
 sky130_fd_sc_hd__and2b_1 _5610_ (.A_N(net2055),
    .B(_2785_),
    .X(_2786_));
 sky130_fd_sc_hd__xor2_1 _5611_ (.A(net2092),
    .B(net2010),
    .X(_2787_));
 sky130_fd_sc_hd__nand2_1 _5612_ (.A(_2786_),
    .B(_2787_),
    .Y(_2788_));
 sky130_fd_sc_hd__nor2_4 _5613_ (.A(net2198),
    .B(_2267_),
    .Y(_2789_));
 sky130_fd_sc_hd__and2_1 _5614_ (.A(net2194),
    .B(_2789_),
    .X(_2790_));
 sky130_fd_sc_hd__nand2_1 _5615_ (.A(net2194),
    .B(_2789_),
    .Y(_2791_));
 sky130_fd_sc_hd__and2_1 _5616_ (.A(net2197),
    .B(_2264_),
    .X(_2792_));
 sky130_fd_sc_hd__nand2_1 _5617_ (.A(net2197),
    .B(_2264_),
    .Y(_2793_));
 sky130_fd_sc_hd__or4b_1 _5618_ (.A(_2785_),
    .B(_2790_),
    .C(_2792_),
    .D_N(_3744_),
    .X(_2794_));
 sky130_fd_sc_hd__a21bo_1 _5619_ (.A1(_2780_),
    .A2(_2784_),
    .B1_N(_2794_),
    .X(_2795_));
 sky130_fd_sc_hd__nand2b_1 _5620_ (.A_N(_2795_),
    .B(_2788_),
    .Y(_2796_));
 sky130_fd_sc_hd__inv_2 _5621_ (.A(_2796_),
    .Y(_2797_));
 sky130_fd_sc_hd__and2_1 _5622_ (.A(net2055),
    .B(_2785_),
    .X(_2798_));
 sky130_fd_sc_hd__nand2_1 _5623_ (.A(net2055),
    .B(_2785_),
    .Y(_2799_));
 sky130_fd_sc_hd__nand2_1 _5624_ (.A(net2092),
    .B(_2798_),
    .Y(_2800_));
 sky130_fd_sc_hd__nor3_1 _5625_ (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .B(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .C(_2791_),
    .Y(_2801_));
 sky130_fd_sc_hd__or3b_1 _5626_ (.A(_2799_),
    .B(net2092),
    .C_N(net2010),
    .X(_2802_));
 sky130_fd_sc_hd__o311a_1 _5627_ (.A1(net2055),
    .A2(net2092),
    .A3(_2791_),
    .B1(_2800_),
    .C1(_2802_),
    .X(_2803_));
 sky130_fd_sc_hd__nand3_1 _5628_ (.A(net2092),
    .B(net2010),
    .C(_2786_),
    .Y(_2804_));
 sky130_fd_sc_hd__o31a_1 _5629_ (.A1(net2092),
    .A2(net2010),
    .A3(_2799_),
    .B1(_2804_),
    .X(_2805_));
 sky130_fd_sc_hd__and3_1 _5630_ (.A(net2240),
    .B(net2234),
    .C(_2789_),
    .X(_2806_));
 sky130_fd_sc_hd__nand2_1 _5631_ (.A(net2055),
    .B(_2790_),
    .Y(_2807_));
 sky130_fd_sc_hd__o2111a_1 _5632_ (.A1(_0068_),
    .A2(_2792_),
    .B1(_2803_),
    .C1(_2805_),
    .D1(_2807_),
    .X(_2808_));
 sky130_fd_sc_hd__and3_1 _5633_ (.A(_2776_),
    .B(_2797_),
    .C(_2808_),
    .X(_0605_));
 sky130_fd_sc_hd__and3_1 _5634_ (.A(_1407_),
    .B(_2776_),
    .C(_2789_),
    .X(_0606_));
 sky130_fd_sc_hd__and3b_1 _5635_ (.A_N(net2197),
    .B(_2776_),
    .C(_2778_),
    .X(_0607_));
 sky130_fd_sc_hd__nand2_4 _5636_ (.A(net2058),
    .B(_2262_),
    .Y(_2809_));
 sky130_fd_sc_hd__nand2_4 _5637_ (.A(net2059),
    .B(_2809_),
    .Y(_2810_));
 sky130_fd_sc_hd__o21ai_1 _5638_ (.A1(_1407_),
    .A2(net2197),
    .B1(net2198),
    .Y(_2811_));
 sky130_fd_sc_hd__o211a_1 _5639_ (.A1(_2267_),
    .A2(_2811_),
    .B1(_2263_),
    .C1(net2059),
    .X(_2812_));
 sky130_fd_sc_hd__nor2_1 _5640_ (.A(net162),
    .B(_2812_),
    .Y(_0608_));
 sky130_fd_sc_hd__and3_1 _5641_ (.A(net801),
    .B(net183),
    .C(net291),
    .X(_0609_));
 sky130_fd_sc_hd__and3_1 _5642_ (.A(net946),
    .B(net181),
    .C(net288),
    .X(_0610_));
 sky130_fd_sc_hd__and3_1 _5643_ (.A(net992),
    .B(net181),
    .C(net288),
    .X(_0611_));
 sky130_fd_sc_hd__and3_1 _5644_ (.A(net894),
    .B(net178),
    .C(net282),
    .X(_0612_));
 sky130_fd_sc_hd__and3_1 _5645_ (.A(net1999),
    .B(net175),
    .C(net278),
    .X(_0613_));
 sky130_fd_sc_hd__and3_1 _5646_ (.A(net944),
    .B(net175),
    .C(net277),
    .X(_0614_));
 sky130_fd_sc_hd__and3_1 _5647_ (.A(net896),
    .B(net178),
    .C(net282),
    .X(_0615_));
 sky130_fd_sc_hd__and3_1 _5648_ (.A(net932),
    .B(net178),
    .C(net282),
    .X(_0616_));
 sky130_fd_sc_hd__and3_1 _5649_ (.A(net902),
    .B(net175),
    .C(net279),
    .X(_0617_));
 sky130_fd_sc_hd__and3_1 _5650_ (.A(net868),
    .B(net175),
    .C(net279),
    .X(_0618_));
 sky130_fd_sc_hd__and3_1 _5651_ (.A(net922),
    .B(net175),
    .C(net277),
    .X(_0619_));
 sky130_fd_sc_hd__and3_1 _5652_ (.A(net974),
    .B(net178),
    .C(net282),
    .X(_0620_));
 sky130_fd_sc_hd__and3_1 _5653_ (.A(net960),
    .B(net178),
    .C(net283),
    .X(_0621_));
 sky130_fd_sc_hd__and3_1 _5654_ (.A(net964),
    .B(net179),
    .C(net285),
    .X(_0622_));
 sky130_fd_sc_hd__and3_1 _5655_ (.A(net2086),
    .B(net2111),
    .C(net287),
    .X(_0623_));
 sky130_fd_sc_hd__and3_1 _5656_ (.A(net1331),
    .B(net2044),
    .C(net285),
    .X(_0624_));
 sky130_fd_sc_hd__and3_1 _5657_ (.A(net713),
    .B(net182),
    .C(net289),
    .X(_0625_));
 sky130_fd_sc_hd__and3_1 _5658_ (.A(net1315),
    .B(net179),
    .C(net286),
    .X(_0626_));
 sky130_fd_sc_hd__and3_1 _5659_ (.A(net906),
    .B(net183),
    .C(net291),
    .X(_0627_));
 sky130_fd_sc_hd__and3_1 _5660_ (.A(net1132),
    .B(net173),
    .C(net276),
    .X(_0628_));
 sky130_fd_sc_hd__and3_1 _5661_ (.A(net942),
    .B(net173),
    .C(net281),
    .X(_0629_));
 sky130_fd_sc_hd__and3_1 _5662_ (.A(net1086),
    .B(net173),
    .C(net276),
    .X(_0630_));
 sky130_fd_sc_hd__and3_1 _5663_ (.A(net870),
    .B(net177),
    .C(net280),
    .X(_0631_));
 sky130_fd_sc_hd__and3_1 _5664_ (.A(net1004),
    .B(net172),
    .C(net274),
    .X(_0632_));
 sky130_fd_sc_hd__and3_1 _5665_ (.A(net1076),
    .B(net172),
    .C(net275),
    .X(_0633_));
 sky130_fd_sc_hd__and3_1 _5666_ (.A(net1108),
    .B(net173),
    .C(net276),
    .X(_0634_));
 sky130_fd_sc_hd__and3_1 _5667_ (.A(net671),
    .B(net171),
    .C(net272),
    .X(_0635_));
 sky130_fd_sc_hd__and3_1 _5668_ (.A(net1028),
    .B(net174),
    .C(net273),
    .X(_0636_));
 sky130_fd_sc_hd__and3_1 _5669_ (.A(net1810),
    .B(net174),
    .C(net273),
    .X(_0637_));
 sky130_fd_sc_hd__and3_1 _5670_ (.A(net1020),
    .B(net173),
    .C(net276),
    .X(_0638_));
 sky130_fd_sc_hd__and3_1 _5671_ (.A(net1357),
    .B(net181),
    .C(net288),
    .X(_0639_));
 sky130_fd_sc_hd__and3_1 _5672_ (.A(net627),
    .B(net181),
    .C(net288),
    .X(_0640_));
 sky130_fd_sc_hd__and3_1 _5673_ (.A(net882),
    .B(net179),
    .C(net284),
    .X(_0641_));
 sky130_fd_sc_hd__and3_1 _5674_ (.A(net978),
    .B(net178),
    .C(net283),
    .X(_0642_));
 sky130_fd_sc_hd__and3_1 _5675_ (.A(net874),
    .B(net175),
    .C(net278),
    .X(_0643_));
 sky130_fd_sc_hd__and3_1 _5676_ (.A(net928),
    .B(net175),
    .C(net277),
    .X(_0644_));
 sky130_fd_sc_hd__and3_1 _5677_ (.A(net643),
    .B(net175),
    .C(net279),
    .X(_0645_));
 sky130_fd_sc_hd__and3_1 _5678_ (.A(net884),
    .B(net179),
    .C(net284),
    .X(_0646_));
 sky130_fd_sc_hd__and3_1 _5679_ (.A(net835),
    .B(net175),
    .C(net279),
    .X(_0647_));
 sky130_fd_sc_hd__and3_1 _5680_ (.A(net845),
    .B(net175),
    .C(net277),
    .X(_0648_));
 sky130_fd_sc_hd__and3_1 _5681_ (.A(net843),
    .B(net178),
    .C(net283),
    .X(_0649_));
 sky130_fd_sc_hd__and3_1 _5682_ (.A(net689),
    .B(net178),
    .C(net283),
    .X(_0650_));
 sky130_fd_sc_hd__and3_1 _5683_ (.A(net1034),
    .B(net179),
    .C(net286),
    .X(_0651_));
 sky130_fd_sc_hd__and3_1 _5684_ (.A(net625),
    .B(net179),
    .C(net285),
    .X(_0652_));
 sky130_fd_sc_hd__and3_1 _5685_ (.A(net701),
    .B(net178),
    .C(net283),
    .X(_0653_));
 sky130_fd_sc_hd__and3_1 _5686_ (.A(net1096),
    .B(net178),
    .C(net284),
    .X(_0654_));
 sky130_fd_sc_hd__and3_1 _5687_ (.A(net880),
    .B(net182),
    .C(net289),
    .X(_0655_));
 sky130_fd_sc_hd__and3_1 _5688_ (.A(net859),
    .B(net180),
    .C(net287),
    .X(_0656_));
 sky130_fd_sc_hd__and3_1 _5689_ (.A(net976),
    .B(net173),
    .C(net274),
    .X(_0657_));
 sky130_fd_sc_hd__and3_1 _5690_ (.A(net956),
    .B(net173),
    .C(net276),
    .X(_0658_));
 sky130_fd_sc_hd__and3_1 _5691_ (.A(net1026),
    .B(net180),
    .C(net287),
    .X(_0659_));
 sky130_fd_sc_hd__and3_1 _5692_ (.A(net912),
    .B(net172),
    .C(net274),
    .X(_0660_));
 sky130_fd_sc_hd__and3_1 _5693_ (.A(net1048),
    .B(net177),
    .C(net280),
    .X(_0661_));
 sky130_fd_sc_hd__and3_1 _5694_ (.A(net1140),
    .B(net172),
    .C(net275),
    .X(_0662_));
 sky130_fd_sc_hd__and3_1 _5695_ (.A(net1208),
    .B(net172),
    .C(net274),
    .X(_0663_));
 sky130_fd_sc_hd__and3_1 _5696_ (.A(net1210),
    .B(net173),
    .C(net276),
    .X(_0664_));
 sky130_fd_sc_hd__and3_1 _5697_ (.A(net926),
    .B(net171),
    .C(net272),
    .X(_0665_));
 sky130_fd_sc_hd__and3_1 _5698_ (.A(net817),
    .B(net171),
    .C(net272),
    .X(_0666_));
 sky130_fd_sc_hd__and3_1 _5699_ (.A(net1170),
    .B(net171),
    .C(net273),
    .X(_0667_));
 sky130_fd_sc_hd__and3_1 _5700_ (.A(net962),
    .B(net177),
    .C(net280),
    .X(_0668_));
 sky130_fd_sc_hd__and3_1 _5701_ (.A(net404),
    .B(net181),
    .C(net290),
    .X(_0669_));
 sky130_fd_sc_hd__and3_1 _5702_ (.A(net397),
    .B(net181),
    .C(net290),
    .X(_0670_));
 sky130_fd_sc_hd__and3_1 _5703_ (.A(net387),
    .B(net181),
    .C(net290),
    .X(_0671_));
 sky130_fd_sc_hd__and3_1 _5704_ (.A(net382),
    .B(net181),
    .C(net290),
    .X(_0672_));
 sky130_fd_sc_hd__and3_1 _5705_ (.A(net433),
    .B(net183),
    .C(net289),
    .X(_0673_));
 sky130_fd_sc_hd__and3_1 _5706_ (.A(net422),
    .B(net2044),
    .C(net289),
    .X(_0674_));
 sky130_fd_sc_hd__and3_1 _5707_ (.A(net414),
    .B(net183),
    .C(net289),
    .X(_0675_));
 sky130_fd_sc_hd__and3_1 _5708_ (.A(net409),
    .B(net182),
    .C(net289),
    .X(_0676_));
 sky130_fd_sc_hd__and3_1 _5709_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[0] ),
    .B(net183),
    .C(net291),
    .X(_0677_));
 sky130_fd_sc_hd__and3_1 _5710_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[1] ),
    .B(net183),
    .C(net291),
    .X(_0678_));
 sky130_fd_sc_hd__and3_1 _5711_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[2] ),
    .B(net183),
    .C(net291),
    .X(_0679_));
 sky130_fd_sc_hd__and3_1 _5712_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[3] ),
    .B(net183),
    .C(net291),
    .X(_0680_));
 sky130_fd_sc_hd__and3_1 _5713_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[4] ),
    .B(net2044),
    .C(net286),
    .X(_0681_));
 sky130_fd_sc_hd__and3_1 _5714_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[5] ),
    .B(net179),
    .C(net285),
    .X(_0682_));
 sky130_fd_sc_hd__and3_1 _5715_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[6] ),
    .B(net177),
    .C(net281),
    .X(_0683_));
 sky130_fd_sc_hd__and3_1 _5716_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[7] ),
    .B(net171),
    .C(net273),
    .X(_0684_));
 sky130_fd_sc_hd__and3_1 _5717_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[8] ),
    .B(net171),
    .C(net273),
    .X(_0685_));
 sky130_fd_sc_hd__and3_1 _5718_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[9] ),
    .B(net2111),
    .C(net287),
    .X(_0686_));
 sky130_fd_sc_hd__and3_1 _5719_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[10] ),
    .B(net175),
    .C(net279),
    .X(_0687_));
 sky130_fd_sc_hd__and3_1 _5720_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[11] ),
    .B(net174),
    .C(net273),
    .X(_0688_));
 sky130_fd_sc_hd__and3_1 _5721_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[12] ),
    .B(net2111),
    .C(net287),
    .X(_0689_));
 sky130_fd_sc_hd__and3_1 _5722_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[13] ),
    .B(net2111),
    .C(net287),
    .X(_0690_));
 sky130_fd_sc_hd__and3_1 _5723_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[14] ),
    .B(net181),
    .C(net290),
    .X(_0691_));
 sky130_fd_sc_hd__and3_1 _5724_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[15] ),
    .B(net179),
    .C(net286),
    .X(_0692_));
 sky130_fd_sc_hd__and3_1 _5725_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[16] ),
    .B(net177),
    .C(net280),
    .X(_0693_));
 sky130_fd_sc_hd__and3_1 _5726_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[17] ),
    .B(net177),
    .C(net281),
    .X(_0694_));
 sky130_fd_sc_hd__and3_1 _5727_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[18] ),
    .B(net181),
    .C(net288),
    .X(_0695_));
 sky130_fd_sc_hd__and3_1 _5728_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[19] ),
    .B(net2111),
    .C(net287),
    .X(_0696_));
 sky130_fd_sc_hd__and3_1 _5729_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[20] ),
    .B(net172),
    .C(net274),
    .X(_0697_));
 sky130_fd_sc_hd__and3_1 _5730_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[21] ),
    .B(net172),
    .C(net275),
    .X(_0698_));
 sky130_fd_sc_hd__and3_1 _5731_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[22] ),
    .B(net183),
    .C(net291),
    .X(_0699_));
 sky130_fd_sc_hd__and3_1 _5732_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[23] ),
    .B(net172),
    .C(net274),
    .X(_0700_));
 sky130_fd_sc_hd__and3_1 _5733_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[24] ),
    .B(net2111),
    .C(net287),
    .X(_0701_));
 sky130_fd_sc_hd__and3_1 _5734_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[25] ),
    .B(net172),
    .C(net274),
    .X(_0702_));
 sky130_fd_sc_hd__and3_1 _5735_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[26] ),
    .B(net172),
    .C(net274),
    .X(_0703_));
 sky130_fd_sc_hd__and3_1 _5736_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[27] ),
    .B(net177),
    .C(net280),
    .X(_0704_));
 sky130_fd_sc_hd__and3_1 _5737_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[28] ),
    .B(net171),
    .C(net273),
    .X(_0705_));
 sky130_fd_sc_hd__and3_1 _5738_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[29] ),
    .B(net171),
    .C(net272),
    .X(_0706_));
 sky130_fd_sc_hd__and3_1 _5739_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[30] ),
    .B(net171),
    .C(net272),
    .X(_0707_));
 sky130_fd_sc_hd__and3_1 _5740_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[31] ),
    .B(net173),
    .C(net276),
    .X(_0708_));
 sky130_fd_sc_hd__and3_1 _5741_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[0] ),
    .B(net183),
    .C(net291),
    .X(_0709_));
 sky130_fd_sc_hd__and3_1 _5742_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[1] ),
    .B(net183),
    .C(net291),
    .X(_0710_));
 sky130_fd_sc_hd__and3_1 _5743_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[2] ),
    .B(net183),
    .C(net291),
    .X(_0711_));
 sky130_fd_sc_hd__and3_1 _5744_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[3] ),
    .B(net181),
    .C(net288),
    .X(_0712_));
 sky130_fd_sc_hd__and3_1 _5745_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[4] ),
    .B(net2111),
    .C(net286),
    .X(_0713_));
 sky130_fd_sc_hd__and3_1 _5746_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[5] ),
    .B(net181),
    .C(net288),
    .X(_0714_));
 sky130_fd_sc_hd__and3_1 _5747_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[6] ),
    .B(net177),
    .C(net281),
    .X(_0715_));
 sky130_fd_sc_hd__and3_1 _5748_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[7] ),
    .B(net171),
    .C(net273),
    .X(_0716_));
 sky130_fd_sc_hd__and3_1 _5749_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[8] ),
    .B(net171),
    .C(net273),
    .X(_0717_));
 sky130_fd_sc_hd__and3_1 _5750_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[9] ),
    .B(net2111),
    .C(net287),
    .X(_0718_));
 sky130_fd_sc_hd__and3_1 _5751_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[10] ),
    .B(net175),
    .C(net279),
    .X(_0719_));
 sky130_fd_sc_hd__and3_1 _5752_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[11] ),
    .B(net174),
    .C(net273),
    .X(_0720_));
 sky130_fd_sc_hd__and3_1 _5753_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[12] ),
    .B(net2111),
    .C(net287),
    .X(_0721_));
 sky130_fd_sc_hd__and3_1 _5754_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[13] ),
    .B(net2111),
    .C(net287),
    .X(_0722_));
 sky130_fd_sc_hd__and3_1 _5755_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[14] ),
    .B(net181),
    .C(net288),
    .X(_0723_));
 sky130_fd_sc_hd__and3_1 _5756_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[15] ),
    .B(net179),
    .C(net286),
    .X(_0724_));
 sky130_fd_sc_hd__and3_1 _5757_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[16] ),
    .B(net177),
    .C(net280),
    .X(_0725_));
 sky130_fd_sc_hd__and3_1 _5758_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[17] ),
    .B(net2111),
    .C(net287),
    .X(_0726_));
 sky130_fd_sc_hd__and3_1 _5759_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[18] ),
    .B(net181),
    .C(net288),
    .X(_0727_));
 sky130_fd_sc_hd__and3_1 _5760_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[19] ),
    .B(net2111),
    .C(net287),
    .X(_0728_));
 sky130_fd_sc_hd__and3_1 _5761_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[20] ),
    .B(net173),
    .C(net274),
    .X(_0729_));
 sky130_fd_sc_hd__and3_1 _5762_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[21] ),
    .B(net172),
    .C(net275),
    .X(_0730_));
 sky130_fd_sc_hd__and3_1 _5763_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[22] ),
    .B(net2111),
    .C(net287),
    .X(_0731_));
 sky130_fd_sc_hd__and3_1 _5764_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[23] ),
    .B(net172),
    .C(net274),
    .X(_0732_));
 sky130_fd_sc_hd__and3_1 _5765_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[24] ),
    .B(net2111),
    .C(net287),
    .X(_0733_));
 sky130_fd_sc_hd__and3_1 _5766_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[25] ),
    .B(net172),
    .C(net274),
    .X(_0734_));
 sky130_fd_sc_hd__and3_1 _5767_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[26] ),
    .B(net172),
    .C(net274),
    .X(_0735_));
 sky130_fd_sc_hd__and3_1 _5768_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[27] ),
    .B(net177),
    .C(net280),
    .X(_0736_));
 sky130_fd_sc_hd__and3_1 _5769_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[28] ),
    .B(net171),
    .C(net272),
    .X(_0737_));
 sky130_fd_sc_hd__and3_1 _5770_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[29] ),
    .B(net171),
    .C(net272),
    .X(_0738_));
 sky130_fd_sc_hd__and3_1 _5771_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[30] ),
    .B(net171),
    .C(net272),
    .X(_0739_));
 sky130_fd_sc_hd__and3_1 _5772_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[31] ),
    .B(net173),
    .C(net276),
    .X(_0740_));
 sky130_fd_sc_hd__and3_1 _5773_ (.A(net2128),
    .B(net182),
    .C(net289),
    .X(_0741_));
 sky130_fd_sc_hd__and3_2 _5774_ (.A(net2204),
    .B(net179),
    .C(net284),
    .X(_0742_));
 sky130_fd_sc_hd__and3_1 _5775_ (.A(net2103),
    .B(net182),
    .C(net290),
    .X(_0743_));
 sky130_fd_sc_hd__and3_1 _5776_ (.A(net2134),
    .B(net182),
    .C(net289),
    .X(_0744_));
 sky130_fd_sc_hd__and3_1 _5777_ (.A(net176),
    .B(net277),
    .C(_2781_),
    .X(_0745_));
 sky130_fd_sc_hd__nor2_1 _5778_ (.A(net162),
    .B(net2195),
    .Y(_0746_));
 sky130_fd_sc_hd__nor2_1 _5779_ (.A(_2263_),
    .B(net162),
    .Y(_0747_));
 sky130_fd_sc_hd__a21o_1 _5780_ (.A1(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ),
    .A2(net2257),
    .B1(net2150),
    .X(_2813_));
 sky130_fd_sc_hd__and3_1 _5781_ (.A(net462),
    .B(net2151),
    .C(net2258),
    .X(_0748_));
 sky130_fd_sc_hd__or2_1 _5782_ (.A(net479),
    .B(_1921_),
    .X(_2814_));
 sky130_fd_sc_hd__a21oi_1 _5783_ (.A1(_1919_),
    .A2(net2151),
    .B1(_2814_),
    .Y(_0749_));
 sky130_fd_sc_hd__and2_1 _5784_ (.A(net469),
    .B(_1931_),
    .X(_0750_));
 sky130_fd_sc_hd__and2_1 _5785_ (.A(net464),
    .B(net2266),
    .X(_0751_));
 sky130_fd_sc_hd__and2_1 _5786_ (.A(net466),
    .B(_1941_),
    .X(_0752_));
 sky130_fd_sc_hd__and2_1 _5787_ (.A(net455),
    .B(_1950_),
    .X(_0753_));
 sky130_fd_sc_hd__and2_1 _5788_ (.A(net456),
    .B(_1959_),
    .X(_0754_));
 sky130_fd_sc_hd__and2_1 _5789_ (.A(net456),
    .B(net2180),
    .X(_0755_));
 sky130_fd_sc_hd__nor2_1 _5790_ (.A(net476),
    .B(net2187),
    .Y(_0756_));
 sky130_fd_sc_hd__and2_1 _5791_ (.A(net456),
    .B(_1988_),
    .X(_0757_));
 sky130_fd_sc_hd__and2_1 _5792_ (.A(net449),
    .B(_1997_),
    .X(_0758_));
 sky130_fd_sc_hd__and2_1 _5793_ (.A(net449),
    .B(_2006_),
    .X(_0759_));
 sky130_fd_sc_hd__and2_1 _5794_ (.A(net455),
    .B(_2015_),
    .X(_0760_));
 sky130_fd_sc_hd__and2_1 _5795_ (.A(net459),
    .B(net2226),
    .X(_0761_));
 sky130_fd_sc_hd__nor2_1 _5796_ (.A(net478),
    .B(_2032_),
    .Y(_0762_));
 sky130_fd_sc_hd__and2_1 _5797_ (.A(net457),
    .B(net2244),
    .X(_0763_));
 sky130_fd_sc_hd__and2_1 _5798_ (.A(net458),
    .B(_2051_),
    .X(_0764_));
 sky130_fd_sc_hd__nor2_1 _5799_ (.A(net478),
    .B(net2255),
    .Y(_0765_));
 sky130_fd_sc_hd__and2_1 _5800_ (.A(net465),
    .B(_2069_),
    .X(_0766_));
 sky130_fd_sc_hd__and2_1 _5801_ (.A(net458),
    .B(net2251),
    .X(_0767_));
 sky130_fd_sc_hd__nor2_1 _5802_ (.A(net480),
    .B(_2087_),
    .Y(_0768_));
 sky130_fd_sc_hd__and2_1 _5803_ (.A(net450),
    .B(net2163),
    .X(_0769_));
 sky130_fd_sc_hd__nor2_1 _5804_ (.A(net474),
    .B(_2106_),
    .Y(_0770_));
 sky130_fd_sc_hd__and2_1 _5805_ (.A(net450),
    .B(net2202),
    .X(_0771_));
 sky130_fd_sc_hd__and2_1 _5806_ (.A(net452),
    .B(_2124_),
    .X(_0772_));
 sky130_fd_sc_hd__and2_1 _5807_ (.A(net445),
    .B(net2126),
    .X(_0773_));
 sky130_fd_sc_hd__and2_1 _5808_ (.A(net445),
    .B(net2219),
    .X(_0774_));
 sky130_fd_sc_hd__and2_1 _5809_ (.A(net450),
    .B(_2151_),
    .X(_0775_));
 sky130_fd_sc_hd__and2_1 _5810_ (.A(net441),
    .B(_2160_),
    .X(_0776_));
 sky130_fd_sc_hd__and2_1 _5811_ (.A(net441),
    .B(net2230),
    .X(_0777_));
 sky130_fd_sc_hd__and2_1 _5812_ (.A(net447),
    .B(net2262),
    .X(_0778_));
 sky130_fd_sc_hd__and2_1 _5813_ (.A(net450),
    .B(net2024),
    .X(_0779_));
 sky130_fd_sc_hd__and2_1 _5814_ (.A(net465),
    .B(net685),
    .X(_0780_));
 sky130_fd_sc_hd__and2_1 _5815_ (.A(net466),
    .B(net681),
    .X(_0781_));
 sky130_fd_sc_hd__and2_1 _5816_ (.A(net465),
    .B(net2027),
    .X(_0782_));
 sky130_fd_sc_hd__and2_1 _5817_ (.A(net465),
    .B(net673),
    .X(_0783_));
 sky130_fd_sc_hd__and2_1 _5818_ (.A(net469),
    .B(net733),
    .X(_0784_));
 sky130_fd_sc_hd__and2_1 _5819_ (.A(net464),
    .B(net775),
    .X(_0785_));
 sky130_fd_sc_hd__and2_1 _5820_ (.A(net464),
    .B(net753),
    .X(_0786_));
 sky130_fd_sc_hd__and2_1 _5821_ (.A(net456),
    .B(net637),
    .X(_0787_));
 sky130_fd_sc_hd__and2_1 _5822_ (.A(net460),
    .B(net853),
    .X(_0788_));
 sky130_fd_sc_hd__and2_1 _5823_ (.A(net456),
    .B(net693),
    .X(_0789_));
 sky130_fd_sc_hd__and2_1 _5824_ (.A(net456),
    .B(net641),
    .X(_0790_));
 sky130_fd_sc_hd__and2_1 _5825_ (.A(net456),
    .B(net749),
    .X(_0791_));
 sky130_fd_sc_hd__and2_1 _5826_ (.A(net449),
    .B(net761),
    .X(_0792_));
 sky130_fd_sc_hd__and2_1 _5827_ (.A(net447),
    .B(net803),
    .X(_0793_));
 sky130_fd_sc_hd__and2_1 _5828_ (.A(net449),
    .B(net747),
    .X(_0794_));
 sky130_fd_sc_hd__and2_1 _5829_ (.A(net456),
    .B(net663),
    .X(_0795_));
 sky130_fd_sc_hd__and2_1 _5830_ (.A(net457),
    .B(net667),
    .X(_0796_));
 sky130_fd_sc_hd__and2_1 _5831_ (.A(net457),
    .B(net649),
    .X(_0797_));
 sky130_fd_sc_hd__and2_1 _5832_ (.A(net462),
    .B(net755),
    .X(_0798_));
 sky130_fd_sc_hd__and2_1 _5833_ (.A(net457),
    .B(net811),
    .X(_0799_));
 sky130_fd_sc_hd__and2_1 _5834_ (.A(net465),
    .B(net727),
    .X(_0800_));
 sky130_fd_sc_hd__and2_1 _5835_ (.A(net458),
    .B(net821),
    .X(_0801_));
 sky130_fd_sc_hd__and2_1 _5836_ (.A(net470),
    .B(net769),
    .X(_0802_));
 sky130_fd_sc_hd__and2_1 _5837_ (.A(net450),
    .B(net793),
    .X(_0803_));
 sky130_fd_sc_hd__and2_1 _5838_ (.A(net451),
    .B(net763),
    .X(_0804_));
 sky130_fd_sc_hd__and2_1 _5839_ (.A(net450),
    .B(net773),
    .X(_0805_));
 sky130_fd_sc_hd__and2_1 _5840_ (.A(net452),
    .B(net743),
    .X(_0806_));
 sky130_fd_sc_hd__and2_1 _5841_ (.A(net445),
    .B(net807),
    .X(_0807_));
 sky130_fd_sc_hd__and2_1 _5842_ (.A(net445),
    .B(net657),
    .X(_0808_));
 sky130_fd_sc_hd__and2_1 _5843_ (.A(net451),
    .B(net886),
    .X(_0809_));
 sky130_fd_sc_hd__and2_1 _5844_ (.A(net441),
    .B(net633),
    .X(_0810_));
 sky130_fd_sc_hd__and2_1 _5845_ (.A(net447),
    .B(net823),
    .X(_0811_));
 sky130_fd_sc_hd__and2_1 _5846_ (.A(net447),
    .B(net699),
    .X(_0812_));
 sky130_fd_sc_hd__and2_1 _5847_ (.A(net451),
    .B(net791),
    .X(_0813_));
 sky130_fd_sc_hd__or3b_4 _5848_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .C_N(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .X(_2815_));
 sky130_fd_sc_hd__nor2_8 _5849_ (.A(_1902_),
    .B(_2815_),
    .Y(_2816_));
 sky130_fd_sc_hd__or2_4 _5850_ (.A(_1902_),
    .B(_2815_),
    .X(_2817_));
 sky130_fd_sc_hd__nor2_2 _5851_ (.A(_1901_),
    .B(_1905_),
    .Y(_2818_));
 sky130_fd_sc_hd__or2_4 _5852_ (.A(_1901_),
    .B(_1905_),
    .X(_2819_));
 sky130_fd_sc_hd__nor2_1 _5853_ (.A(_2816_),
    .B(_2818_),
    .Y(_2820_));
 sky130_fd_sc_hd__nand2_4 _5854_ (.A(_2817_),
    .B(_2819_),
    .Y(_2821_));
 sky130_fd_sc_hd__mux4_1 _5855_ (.A0(_1674_),
    .A1(_1701_),
    .A2(_1662_),
    .A3(_1689_),
    .S0(net201),
    .S1(net196),
    .X(_2822_));
 sky130_fd_sc_hd__mux4_1 _5856_ (.A0(_1723_),
    .A1(_1733_),
    .A2(_1749_),
    .A3(_1712_),
    .S0(net199),
    .S1(net195),
    .X(_2823_));
 sky130_fd_sc_hd__or2_1 _5857_ (.A(net204),
    .B(_2822_),
    .X(_2824_));
 sky130_fd_sc_hd__o211a_1 _5858_ (.A1(net207),
    .A2(_2823_),
    .B1(_2824_),
    .C1(net214),
    .X(_2825_));
 sky130_fd_sc_hd__mux2_1 _5859_ (.A0(_1772_),
    .A1(_1793_),
    .S(net193),
    .X(_2826_));
 sky130_fd_sc_hd__mux4_1 _5860_ (.A0(_1772_),
    .A1(_1793_),
    .A2(_1783_),
    .A3(_1762_),
    .S0(net195),
    .S1(net200),
    .X(_2827_));
 sky130_fd_sc_hd__mux2_1 _5861_ (.A0(_1828_),
    .A1(_1806_),
    .S(net193),
    .X(_2828_));
 sky130_fd_sc_hd__mux2_1 _5862_ (.A0(_1815_),
    .A1(_1839_),
    .S(net193),
    .X(_2829_));
 sky130_fd_sc_hd__mux2_1 _5863_ (.A0(_2828_),
    .A1(_2829_),
    .S(net198),
    .X(_2830_));
 sky130_fd_sc_hd__mux2_1 _5864_ (.A0(_2827_),
    .A1(_2830_),
    .S(net203),
    .X(_2831_));
 sky130_fd_sc_hd__mux2_1 _5865_ (.A0(_1544_),
    .A1(_1521_),
    .S(net194),
    .X(_2832_));
 sky130_fd_sc_hd__mux2_1 _5866_ (.A0(_1555_),
    .A1(_1531_),
    .S(net193),
    .X(_2833_));
 sky130_fd_sc_hd__mux2_1 _5867_ (.A0(_2832_),
    .A1(_2833_),
    .S(net198),
    .X(_2834_));
 sky130_fd_sc_hd__mux2_1 _5868_ (.A0(_1590_),
    .A1(_1567_),
    .S(net193),
    .X(_2835_));
 sky130_fd_sc_hd__mux2_1 _5869_ (.A0(_1577_),
    .A1(_1601_),
    .S(net192),
    .X(_2836_));
 sky130_fd_sc_hd__mux2_1 _5870_ (.A0(_2835_),
    .A1(_2836_),
    .S(net197),
    .X(_2837_));
 sky130_fd_sc_hd__mux2_1 _5871_ (.A0(_2834_),
    .A1(_2837_),
    .S(net203),
    .X(_2838_));
 sky130_fd_sc_hd__mux2_1 _5872_ (.A0(_1637_),
    .A1(_1614_),
    .S(net192),
    .X(_2839_));
 sky130_fd_sc_hd__mux2_1 _5873_ (.A0(_1624_),
    .A1(_1649_),
    .S(net192),
    .X(_2840_));
 sky130_fd_sc_hd__mux2_1 _5874_ (.A0(_2839_),
    .A1(_2840_),
    .S(net197),
    .X(_2841_));
 sky130_fd_sc_hd__mux2_1 _5875_ (.A0(_1480_),
    .A1(_1503_),
    .S(net192),
    .X(_2842_));
 sky130_fd_sc_hd__mux2_1 _5876_ (.A0(_1490_),
    .A1(_1467_),
    .S(net192),
    .X(_2843_));
 sky130_fd_sc_hd__mux2_1 _5877_ (.A0(_2842_),
    .A1(_2843_),
    .S(net197),
    .X(_2844_));
 sky130_fd_sc_hd__mux2_1 _5878_ (.A0(_2841_),
    .A1(_2844_),
    .S(net202),
    .X(_2845_));
 sky130_fd_sc_hd__mux2_2 _5879_ (.A0(_2838_),
    .A1(_2845_),
    .S(net209),
    .X(_2846_));
 sky130_fd_sc_hd__a211o_1 _5880_ (.A1(net210),
    .A2(_2831_),
    .B1(_2825_),
    .C1(net187),
    .X(_2847_));
 sky130_fd_sc_hd__o211ai_2 _5881_ (.A1(net191),
    .A2(_2846_),
    .B1(_2847_),
    .C1(_2821_),
    .Y(_2848_));
 sky130_fd_sc_hd__or3_1 _5882_ (.A(net210),
    .B(net204),
    .C(_1852_),
    .X(_2849_));
 sky130_fd_sc_hd__nor2_8 _5883_ (.A(_1901_),
    .B(_2815_),
    .Y(_2850_));
 sky130_fd_sc_hd__or2_4 _5884_ (.A(_1901_),
    .B(_2815_),
    .X(_2851_));
 sky130_fd_sc_hd__nor2_1 _5885_ (.A(net187),
    .B(_2851_),
    .Y(_2852_));
 sky130_fd_sc_hd__nand2_4 _5886_ (.A(net190),
    .B(_2850_),
    .Y(_2853_));
 sky130_fd_sc_hd__nor2_1 _5887_ (.A(net2188),
    .B(net2346),
    .Y(_2854_));
 sky130_fd_sc_hd__or2_2 _5888_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .X(_2855_));
 sky130_fd_sc_hd__nor2_2 _5889_ (.A(_2815_),
    .B(_2855_),
    .Y(_2856_));
 sky130_fd_sc_hd__and4bb_2 _5890_ (.A_N(net2293),
    .B_N(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .C(net2232),
    .D(_2854_),
    .X(_2857_));
 sky130_fd_sc_hd__or4_1 _5891_ (.A(_2821_),
    .B(_2850_),
    .C(net364),
    .D(net362),
    .X(_2858_));
 sky130_fd_sc_hd__nor2_8 _5892_ (.A(_1901_),
    .B(_1903_),
    .Y(_2859_));
 sky130_fd_sc_hd__or2_1 _5893_ (.A(_1901_),
    .B(_1903_),
    .X(_2860_));
 sky130_fd_sc_hd__a21oi_4 _5894_ (.A1(_1899_),
    .A2(_2854_),
    .B1(_2859_),
    .Y(_2861_));
 sky130_fd_sc_hd__inv_4 _5895_ (.A(net319),
    .Y(_2862_));
 sky130_fd_sc_hd__nor2_4 _5896_ (.A(_1905_),
    .B(_2855_),
    .Y(_2863_));
 sky130_fd_sc_hd__or2_4 _5897_ (.A(_1905_),
    .B(_2855_),
    .X(_2864_));
 sky130_fd_sc_hd__nand2_1 _5898_ (.A(net319),
    .B(_2864_),
    .Y(_2865_));
 sky130_fd_sc_hd__and4b_1 _5899_ (.A_N(_2858_),
    .B(_2864_),
    .C(net319),
    .D(_1906_),
    .X(_2866_));
 sky130_fd_sc_hd__or4b_2 _5900_ (.A(_2858_),
    .B(net358),
    .C(_2862_),
    .D_N(_1906_),
    .X(_2867_));
 sky130_fd_sc_hd__a221o_1 _5901_ (.A1(net196),
    .A2(net362),
    .B1(_2865_),
    .B2(_1703_),
    .C1(net364),
    .X(_2868_));
 sky130_fd_sc_hd__a21oi_1 _5902_ (.A1(_1704_),
    .A2(_2868_),
    .B1(net224),
    .Y(_2869_));
 sky130_fd_sc_hd__o221a_1 _5903_ (.A1(_1896_),
    .A2(_1904_),
    .B1(_2849_),
    .B2(_2853_),
    .C1(_2869_),
    .X(_2870_));
 sky130_fd_sc_hd__a221oi_2 _5904_ (.A1(_1703_),
    .A2(net224),
    .B1(net2355),
    .B2(_2848_),
    .C1(net476),
    .Y(_0814_));
 sky130_fd_sc_hd__mux4_1 _5905_ (.A0(_1567_),
    .A1(_1577_),
    .A2(_1601_),
    .A3(_1637_),
    .S0(net192),
    .S1(net197),
    .X(_2871_));
 sky130_fd_sc_hd__mux2_1 _5906_ (.A0(_1521_),
    .A1(_1555_),
    .S(net193),
    .X(_2872_));
 sky130_fd_sc_hd__mux4_1 _5907_ (.A0(_1521_),
    .A1(_1531_),
    .A2(_1555_),
    .A3(_1590_),
    .S0(net198),
    .S1(net193),
    .X(_2873_));
 sky130_fd_sc_hd__mux2_1 _5908_ (.A0(_2871_),
    .A1(_2873_),
    .S(net206),
    .X(_2874_));
 sky130_fd_sc_hd__nor2_1 _5909_ (.A(net209),
    .B(_2874_),
    .Y(_2875_));
 sky130_fd_sc_hd__mux4_1 _5910_ (.A0(_1614_),
    .A1(_1624_),
    .A2(_1649_),
    .A3(_1480_),
    .S0(net194),
    .S1(net197),
    .X(_2876_));
 sky130_fd_sc_hd__nor2_1 _5911_ (.A(net202),
    .B(_2876_),
    .Y(_2877_));
 sky130_fd_sc_hd__mux2_1 _5912_ (.A0(_1503_),
    .A1(_1490_),
    .S(net194),
    .X(_2878_));
 sky130_fd_sc_hd__and2_1 _5913_ (.A(net200),
    .B(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__a21oi_1 _5914_ (.A1(_1467_),
    .A2(net197),
    .B1(_2879_),
    .Y(_2880_));
 sky130_fd_sc_hd__a21o_1 _5915_ (.A1(net202),
    .A2(_2880_),
    .B1(_2877_),
    .X(_2881_));
 sky130_fd_sc_hd__a21oi_1 _5916_ (.A1(net209),
    .A2(_2881_),
    .B1(_2875_),
    .Y(_2882_));
 sky130_fd_sc_hd__a31oi_2 _5917_ (.A1(_1467_),
    .A2(net197),
    .A3(_1699_),
    .B1(_2879_),
    .Y(_2883_));
 sky130_fd_sc_hd__a21oi_2 _5918_ (.A1(net202),
    .A2(_2883_),
    .B1(_2877_),
    .Y(_2884_));
 sky130_fd_sc_hd__o21ba_1 _5919_ (.A1(net213),
    .A2(_2884_),
    .B1_N(_2875_),
    .X(_2885_));
 sky130_fd_sc_hd__a22o_1 _5920_ (.A1(_2816_),
    .A2(_2882_),
    .B1(_2885_),
    .B2(_2818_),
    .X(_2886_));
 sky130_fd_sc_hd__or3_1 _5921_ (.A(_1683_),
    .B(_1685_),
    .C(_2859_),
    .X(_2887_));
 sky130_fd_sc_hd__o21ai_1 _5922_ (.A1(_1683_),
    .A2(_1685_),
    .B1(_2859_),
    .Y(_2888_));
 sky130_fd_sc_hd__and3_1 _5923_ (.A(_1689_),
    .B(_2887_),
    .C(_2888_),
    .X(_2889_));
 sky130_fd_sc_hd__a21o_1 _5924_ (.A1(_2887_),
    .A2(_2888_),
    .B1(_1689_),
    .X(_2890_));
 sky130_fd_sc_hd__and2b_1 _5925_ (.A_N(_2889_),
    .B(_2890_),
    .X(_2891_));
 sky130_fd_sc_hd__mux2_1 _5926_ (.A0(_2859_),
    .A1(_1701_),
    .S(net196),
    .X(_2892_));
 sky130_fd_sc_hd__xor2_1 _5927_ (.A(_2891_),
    .B(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__a221o_1 _5928_ (.A1(_1691_),
    .A2(net364),
    .B1(net362),
    .B2(net199),
    .C1(net224),
    .X(_2894_));
 sky130_fd_sc_hd__mux2_1 _5929_ (.A0(_1689_),
    .A1(_1701_),
    .S(net196),
    .X(_2895_));
 sky130_fd_sc_hd__nand2_1 _5930_ (.A(net201),
    .B(_2895_),
    .Y(_2896_));
 sky130_fd_sc_hd__or2_1 _5931_ (.A(net204),
    .B(_2896_),
    .X(_2897_));
 sky130_fd_sc_hd__or2_1 _5932_ (.A(net210),
    .B(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__a2bb2o_1 _5933_ (.A1_N(_2853_),
    .A2_N(_2898_),
    .B1(_2893_),
    .B2(_2862_),
    .X(_2899_));
 sky130_fd_sc_hd__a211o_1 _5934_ (.A1(net358),
    .A2(_2891_),
    .B1(_2894_),
    .C1(_2899_),
    .X(_2900_));
 sky130_fd_sc_hd__mux4_1 _5935_ (.A0(_1662_),
    .A1(_1689_),
    .A2(_1723_),
    .A3(_1674_),
    .S0(net201),
    .S1(net196),
    .X(_2901_));
 sky130_fd_sc_hd__mux4_1 _5936_ (.A0(_1712_),
    .A1(_1749_),
    .A2(_1783_),
    .A3(_1733_),
    .S0(net201),
    .S1(net195),
    .X(_2902_));
 sky130_fd_sc_hd__mux2_1 _5937_ (.A0(_2901_),
    .A1(_2902_),
    .S(net204),
    .X(_2903_));
 sky130_fd_sc_hd__mux2_1 _5938_ (.A0(_1806_),
    .A1(_1815_),
    .S(net194),
    .X(_2904_));
 sky130_fd_sc_hd__mux2_1 _5939_ (.A0(_1839_),
    .A1(_1544_),
    .S(net193),
    .X(_2905_));
 sky130_fd_sc_hd__mux2_1 _5940_ (.A0(_2904_),
    .A1(_2905_),
    .S(net198),
    .X(_2906_));
 sky130_fd_sc_hd__mux2_1 _5941_ (.A0(_1793_),
    .A1(_1828_),
    .S(net194),
    .X(_2907_));
 sky130_fd_sc_hd__mux4_1 _5942_ (.A0(_1762_),
    .A1(_1772_),
    .A2(_1793_),
    .A3(_1828_),
    .S0(net195),
    .S1(net198),
    .X(_2908_));
 sky130_fd_sc_hd__mux2_1 _5943_ (.A0(_2906_),
    .A1(_2908_),
    .S(net206),
    .X(_2909_));
 sky130_fd_sc_hd__mux2_1 _5944_ (.A0(_2903_),
    .A1(_2909_),
    .S(net211),
    .X(_2910_));
 sky130_fd_sc_hd__nor2_1 _5945_ (.A(net188),
    .B(_2820_),
    .Y(_2911_));
 sky130_fd_sc_hd__a221o_1 _5946_ (.A1(net188),
    .A2(_2886_),
    .B1(_2910_),
    .B2(_2911_),
    .C1(_2900_),
    .X(_2912_));
 sky130_fd_sc_hd__a21o_1 _5947_ (.A1(net199),
    .A2(_1689_),
    .B1(net222),
    .X(_2913_));
 sky130_fd_sc_hd__and3_1 _5948_ (.A(net461),
    .B(_2912_),
    .C(_2913_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_1 _5949_ (.A0(_1674_),
    .A1(_1689_),
    .S(net196),
    .X(_2914_));
 sky130_fd_sc_hd__o21bai_1 _5950_ (.A1(net199),
    .A2(_2914_),
    .B1_N(_1851_),
    .Y(_2915_));
 sky130_fd_sc_hd__nor2_1 _5951_ (.A(net204),
    .B(_2915_),
    .Y(_2916_));
 sky130_fd_sc_hd__mux4_1 _5952_ (.A0(_1674_),
    .A1(_1723_),
    .A2(_1662_),
    .A3(_1749_),
    .S0(net199),
    .S1(net195),
    .X(_2917_));
 sky130_fd_sc_hd__mux4_1 _5953_ (.A0(_1733_),
    .A1(_1783_),
    .A2(_1712_),
    .A3(_1762_),
    .S0(net199),
    .S1(net195),
    .X(_2918_));
 sky130_fd_sc_hd__mux2_1 _5954_ (.A0(_2917_),
    .A1(_2918_),
    .S(net204),
    .X(_2919_));
 sky130_fd_sc_hd__mux2_1 _5955_ (.A0(_2826_),
    .A1(_2828_),
    .S(net198),
    .X(_2920_));
 sky130_fd_sc_hd__mux2_1 _5956_ (.A0(_2829_),
    .A1(_2832_),
    .S(net198),
    .X(_2921_));
 sky130_fd_sc_hd__mux2_1 _5957_ (.A0(_2920_),
    .A1(_2921_),
    .S(net203),
    .X(_2922_));
 sky130_fd_sc_hd__mux2_1 _5958_ (.A0(_2919_),
    .A1(_2922_),
    .S(net210),
    .X(_2923_));
 sky130_fd_sc_hd__a32o_1 _5959_ (.A1(net214),
    .A2(_2850_),
    .A3(_2916_),
    .B1(_2923_),
    .B2(_2821_),
    .X(_2924_));
 sky130_fd_sc_hd__nand2_1 _5960_ (.A(net191),
    .B(_2924_),
    .Y(_2925_));
 sky130_fd_sc_hd__mux2_1 _5961_ (.A0(_2840_),
    .A1(_2842_),
    .S(net197),
    .X(_2926_));
 sky130_fd_sc_hd__or2_1 _5962_ (.A(net202),
    .B(_2926_),
    .X(_2927_));
 sky130_fd_sc_hd__nand2_1 _5963_ (.A(net200),
    .B(_2843_),
    .Y(_2928_));
 sky130_fd_sc_hd__a21boi_2 _5964_ (.A1(net202),
    .A2(_2928_),
    .B1_N(_2927_),
    .Y(_2929_));
 sky130_fd_sc_hd__inv_2 _5965_ (.A(_2929_),
    .Y(_2930_));
 sky130_fd_sc_hd__mux2_1 _5966_ (.A0(_2833_),
    .A1(_2835_),
    .S(net198),
    .X(_2931_));
 sky130_fd_sc_hd__mux2_1 _5967_ (.A0(_2836_),
    .A1(_2839_),
    .S(net197),
    .X(_2932_));
 sky130_fd_sc_hd__mux2_1 _5968_ (.A0(_2931_),
    .A1(_2932_),
    .S(net203),
    .X(_2933_));
 sky130_fd_sc_hd__nor2_1 _5969_ (.A(net209),
    .B(_2933_),
    .Y(_2934_));
 sky130_fd_sc_hd__a211o_1 _5970_ (.A1(net209),
    .A2(_2930_),
    .B1(_2934_),
    .C1(_2819_),
    .X(_2935_));
 sky130_fd_sc_hd__o21ai_1 _5971_ (.A1(_1468_),
    .A2(net200),
    .B1(_2928_),
    .Y(_2936_));
 sky130_fd_sc_hd__o21ai_1 _5972_ (.A1(net205),
    .A2(_2936_),
    .B1(_2927_),
    .Y(_2937_));
 sky130_fd_sc_hd__a211o_1 _5973_ (.A1(net209),
    .A2(_2937_),
    .B1(_2934_),
    .C1(_2817_),
    .X(_2938_));
 sky130_fd_sc_hd__a21o_1 _5974_ (.A1(_2935_),
    .A2(_2938_),
    .B1(net190),
    .X(_2939_));
 sky130_fd_sc_hd__o21a_1 _5975_ (.A1(_2889_),
    .A2(_2892_),
    .B1(_2890_),
    .X(_2940_));
 sky130_fd_sc_hd__nand2_1 _5976_ (.A(net207),
    .B(net360),
    .Y(_2941_));
 sky130_fd_sc_hd__nand2_1 _5977_ (.A(net204),
    .B(_2859_),
    .Y(_2942_));
 sky130_fd_sc_hd__and3_1 _5978_ (.A(_1674_),
    .B(_2941_),
    .C(_2942_),
    .X(_2943_));
 sky130_fd_sc_hd__a21o_1 _5979_ (.A1(_2941_),
    .A2(_2942_),
    .B1(_1674_),
    .X(_2944_));
 sky130_fd_sc_hd__and2b_1 _5980_ (.A_N(_2943_),
    .B(_2944_),
    .X(_2945_));
 sky130_fd_sc_hd__xnor2_1 _5981_ (.A(_2940_),
    .B(_2945_),
    .Y(_2946_));
 sky130_fd_sc_hd__a221o_1 _5982_ (.A1(net204),
    .A2(_2857_),
    .B1(_2863_),
    .B2(_1675_),
    .C1(_2856_),
    .X(_2947_));
 sky130_fd_sc_hd__o21ai_1 _5983_ (.A1(net204),
    .A2(_1674_),
    .B1(_2947_),
    .Y(_2948_));
 sky130_fd_sc_hd__o2111a_1 _5984_ (.A1(net319),
    .A2(_2946_),
    .B1(_2948_),
    .C1(net222),
    .D1(_2939_),
    .X(_2949_));
 sky130_fd_sc_hd__a221oi_2 _5985_ (.A1(net2334),
    .A2(net225),
    .B1(_2925_),
    .B2(_2949_),
    .C1(net479),
    .Y(_0816_));
 sky130_fd_sc_hd__mux4_1 _5986_ (.A0(_1531_),
    .A1(_1567_),
    .A2(_1590_),
    .A3(_1577_),
    .S0(net198),
    .S1(net193),
    .X(_2950_));
 sky130_fd_sc_hd__mux4_1 _5987_ (.A0(_1601_),
    .A1(_1614_),
    .A2(_1637_),
    .A3(_1624_),
    .S0(net197),
    .S1(net192),
    .X(_2951_));
 sky130_fd_sc_hd__mux2_1 _5988_ (.A0(_2950_),
    .A1(_2951_),
    .S(net202),
    .X(_2952_));
 sky130_fd_sc_hd__mux4_1 _5989_ (.A0(_1649_),
    .A1(_1503_),
    .A2(_1480_),
    .A3(_1490_),
    .S0(net197),
    .S1(net192),
    .X(_2953_));
 sky130_fd_sc_hd__nand2_1 _5990_ (.A(net205),
    .B(_2953_),
    .Y(_2954_));
 sky130_fd_sc_hd__nand2_1 _5991_ (.A(_1467_),
    .B(net202),
    .Y(_2955_));
 sky130_fd_sc_hd__nand2_1 _5992_ (.A(_2954_),
    .B(_2955_),
    .Y(_2956_));
 sky130_fd_sc_hd__mux2_1 _5993_ (.A0(_2952_),
    .A1(_2956_),
    .S(net208),
    .X(_2957_));
 sky130_fd_sc_hd__or3_1 _5994_ (.A(_1468_),
    .B(net197),
    .C(net192),
    .X(_2958_));
 sky130_fd_sc_hd__o21a_1 _5995_ (.A1(net205),
    .A2(_2958_),
    .B1(_2954_),
    .X(_2959_));
 sky130_fd_sc_hd__inv_2 _5996_ (.A(_2959_),
    .Y(_2960_));
 sky130_fd_sc_hd__mux2_1 _5997_ (.A0(_2952_),
    .A1(_2960_),
    .S(net208),
    .X(_2961_));
 sky130_fd_sc_hd__a22o_1 _5998_ (.A1(_2816_),
    .A2(_2957_),
    .B1(_2961_),
    .B2(_2818_),
    .X(_2962_));
 sky130_fd_sc_hd__xnor2_1 _5999_ (.A(_1659_),
    .B(_2859_),
    .Y(_2963_));
 sky130_fd_sc_hd__and2_1 _6000_ (.A(_1662_),
    .B(_2963_),
    .X(_2964_));
 sky130_fd_sc_hd__or2_1 _6001_ (.A(_1662_),
    .B(_2963_),
    .X(_2965_));
 sky130_fd_sc_hd__and2b_1 _6002_ (.A_N(_2964_),
    .B(_2965_),
    .X(_2966_));
 sky130_fd_sc_hd__o21a_1 _6003_ (.A1(_2940_),
    .A2(_2943_),
    .B1(_2944_),
    .X(_2967_));
 sky130_fd_sc_hd__xnor2_1 _6004_ (.A(_2966_),
    .B(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__nor2_1 _6005_ (.A(_2861_),
    .B(_2968_),
    .Y(_2969_));
 sky130_fd_sc_hd__mux2_1 _6006_ (.A0(_1662_),
    .A1(_1674_),
    .S(net196),
    .X(_2970_));
 sky130_fd_sc_hd__mux2_1 _6007_ (.A0(_2895_),
    .A1(_2970_),
    .S(net201),
    .X(_2971_));
 sky130_fd_sc_hd__nand2_1 _6008_ (.A(net207),
    .B(_2971_),
    .Y(_2972_));
 sky130_fd_sc_hd__or2_1 _6009_ (.A(net210),
    .B(_2972_),
    .X(_2973_));
 sky130_fd_sc_hd__nor2_1 _6010_ (.A(_2853_),
    .B(_2973_),
    .Y(_2974_));
 sky130_fd_sc_hd__a221o_1 _6011_ (.A1(_1663_),
    .A2(net364),
    .B1(net362),
    .B2(net211),
    .C1(net225),
    .X(_2975_));
 sky130_fd_sc_hd__a21o_1 _6012_ (.A1(_2863_),
    .A2(_2966_),
    .B1(_2975_),
    .X(_2976_));
 sky130_fd_sc_hd__mux4_1 _6013_ (.A0(_1662_),
    .A1(_1723_),
    .A2(_1749_),
    .A3(_1733_),
    .S0(net196),
    .S1(net199),
    .X(_2977_));
 sky130_fd_sc_hd__mux4_1 _6014_ (.A0(_1712_),
    .A1(_1762_),
    .A2(_1783_),
    .A3(_1772_),
    .S0(net198),
    .S1(net193),
    .X(_2978_));
 sky130_fd_sc_hd__mux2_1 _6015_ (.A0(_2977_),
    .A1(_2978_),
    .S(net204),
    .X(_2979_));
 sky130_fd_sc_hd__mux2_1 _6016_ (.A0(_2904_),
    .A1(_2907_),
    .S(net200),
    .X(_2980_));
 sky130_fd_sc_hd__mux2_1 _6017_ (.A0(_2872_),
    .A1(_2905_),
    .S(net200),
    .X(_2981_));
 sky130_fd_sc_hd__mux2_1 _6018_ (.A0(_2980_),
    .A1(_2981_),
    .S(net203),
    .X(_2982_));
 sky130_fd_sc_hd__mux2_1 _6019_ (.A0(_2979_),
    .A1(_2982_),
    .S(net210),
    .X(_2983_));
 sky130_fd_sc_hd__a211o_1 _6020_ (.A1(_2911_),
    .A2(_2983_),
    .B1(_2976_),
    .C1(_2974_),
    .X(_2984_));
 sky130_fd_sc_hd__a211o_1 _6021_ (.A1(net188),
    .A2(_2962_),
    .B1(_2969_),
    .C1(_2984_),
    .X(_2985_));
 sky130_fd_sc_hd__a21o_1 _6022_ (.A1(net211),
    .A2(_1662_),
    .B1(net222),
    .X(_2986_));
 sky130_fd_sc_hd__and3_1 _6023_ (.A(net461),
    .B(_2985_),
    .C(_2986_),
    .X(_0817_));
 sky130_fd_sc_hd__o21ai_2 _6024_ (.A1(_2964_),
    .A2(_2967_),
    .B1(_2965_),
    .Y(_2987_));
 sky130_fd_sc_hd__xnor2_1 _6025_ (.A(net191),
    .B(_2859_),
    .Y(_2988_));
 sky130_fd_sc_hd__nand2_1 _6026_ (.A(_1723_),
    .B(_2988_),
    .Y(_2989_));
 sky130_fd_sc_hd__nor2_1 _6027_ (.A(_1723_),
    .B(_2988_),
    .Y(_2990_));
 sky130_fd_sc_hd__or2_1 _6028_ (.A(_1723_),
    .B(_2988_),
    .X(_2991_));
 sky130_fd_sc_hd__nand2_1 _6029_ (.A(_2989_),
    .B(_2991_),
    .Y(_2992_));
 sky130_fd_sc_hd__and2_1 _6030_ (.A(_2987_),
    .B(_2992_),
    .X(_2993_));
 sky130_fd_sc_hd__nor2_1 _6031_ (.A(_2987_),
    .B(_2992_),
    .Y(_2994_));
 sky130_fd_sc_hd__mux2_1 _6032_ (.A0(_2837_),
    .A1(_2841_),
    .S(net202),
    .X(_2995_));
 sky130_fd_sc_hd__and2_1 _6033_ (.A(net205),
    .B(_2844_),
    .X(_2996_));
 sky130_fd_sc_hd__a21oi_1 _6034_ (.A1(_1467_),
    .A2(net202),
    .B1(_2996_),
    .Y(_2997_));
 sky130_fd_sc_hd__inv_2 _6035_ (.A(_2997_),
    .Y(_2998_));
 sky130_fd_sc_hd__mux2_1 _6036_ (.A0(_2995_),
    .A1(_2998_),
    .S(net208),
    .X(_2999_));
 sky130_fd_sc_hd__o311a_1 _6037_ (.A1(net212),
    .A2(_2816_),
    .A3(_2996_),
    .B1(_2999_),
    .C1(net185),
    .X(_3000_));
 sky130_fd_sc_hd__mux2_1 _6038_ (.A0(_2830_),
    .A1(_2834_),
    .S(net203),
    .X(_3001_));
 sky130_fd_sc_hd__mux2_1 _6039_ (.A0(_2823_),
    .A1(_2827_),
    .S(net204),
    .X(_3002_));
 sky130_fd_sc_hd__or2_1 _6040_ (.A(net209),
    .B(_3002_),
    .X(_3003_));
 sky130_fd_sc_hd__o211a_1 _6041_ (.A1(net214),
    .A2(_3001_),
    .B1(_3003_),
    .C1(net191),
    .X(_3004_));
 sky130_fd_sc_hd__o21ai_1 _6042_ (.A1(_3000_),
    .A2(_3004_),
    .B1(_2821_),
    .Y(_3005_));
 sky130_fd_sc_hd__mux4_1 _6043_ (.A0(_1674_),
    .A1(_1723_),
    .A2(_1689_),
    .A3(_1662_),
    .S0(net201),
    .S1(net196),
    .X(_3006_));
 sky130_fd_sc_hd__nor2_1 _6044_ (.A(net204),
    .B(_3006_),
    .Y(_3007_));
 sky130_fd_sc_hd__a21o_1 _6045_ (.A1(net204),
    .A2(_1852_),
    .B1(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__or2_1 _6046_ (.A(net211),
    .B(_3008_),
    .X(_3009_));
 sky130_fd_sc_hd__a221o_1 _6047_ (.A1(net188),
    .A2(net362),
    .B1(net358),
    .B2(_1724_),
    .C1(net364),
    .X(_3010_));
 sky130_fd_sc_hd__nand2_1 _6048_ (.A(_1725_),
    .B(_3010_),
    .Y(_3011_));
 sky130_fd_sc_hd__o211a_1 _6049_ (.A1(_2853_),
    .A2(_3009_),
    .B1(_3011_),
    .C1(net222),
    .X(_3012_));
 sky130_fd_sc_hd__o311a_1 _6050_ (.A1(net2347),
    .A2(_2993_),
    .A3(_2994_),
    .B1(_3005_),
    .C1(_3012_),
    .X(_3013_));
 sky130_fd_sc_hd__a211oi_1 _6051_ (.A1(_1724_),
    .A2(net224),
    .B1(_3013_),
    .C1(net476),
    .Y(_0818_));
 sky130_fd_sc_hd__xnor2_1 _6052_ (.A(_1747_),
    .B(net360),
    .Y(_3014_));
 sky130_fd_sc_hd__nor2_1 _6053_ (.A(_1749_),
    .B(_3014_),
    .Y(_3015_));
 sky130_fd_sc_hd__nand2_1 _6054_ (.A(_1749_),
    .B(_3014_),
    .Y(_3016_));
 sky130_fd_sc_hd__nand2b_1 _6055_ (.A_N(_3015_),
    .B(_3016_),
    .Y(_3017_));
 sky130_fd_sc_hd__a21o_1 _6056_ (.A1(_2987_),
    .A2(_2989_),
    .B1(_2990_),
    .X(_3018_));
 sky130_fd_sc_hd__xnor2_1 _6057_ (.A(_3017_),
    .B(_3018_),
    .Y(_3019_));
 sky130_fd_sc_hd__mux2_1 _6058_ (.A0(_2871_),
    .A1(_2876_),
    .S(net202),
    .X(_3020_));
 sky130_fd_sc_hd__nor2_1 _6059_ (.A(net208),
    .B(_3020_),
    .Y(_3021_));
 sky130_fd_sc_hd__o21a_1 _6060_ (.A1(net202),
    .A2(_2880_),
    .B1(_2955_),
    .X(_3022_));
 sky130_fd_sc_hd__a21o_1 _6061_ (.A1(net208),
    .A2(_3022_),
    .B1(_3021_),
    .X(_3023_));
 sky130_fd_sc_hd__nor2_1 _6062_ (.A(_2817_),
    .B(_3023_),
    .Y(_3024_));
 sky130_fd_sc_hd__or2_2 _6063_ (.A(net202),
    .B(_2883_),
    .X(_3025_));
 sky130_fd_sc_hd__a211oi_4 _6064_ (.A1(net208),
    .A2(_3025_),
    .B1(_3021_),
    .C1(_2819_),
    .Y(_3026_));
 sky130_fd_sc_hd__o21ai_4 _6065_ (.A1(_3024_),
    .A2(_3026_),
    .B1(net185),
    .Y(_3027_));
 sky130_fd_sc_hd__a221oi_1 _6066_ (.A1(_1750_),
    .A2(net364),
    .B1(net362),
    .B2(_1747_),
    .C1(net224),
    .Y(_3028_));
 sky130_fd_sc_hd__mux2_1 _6067_ (.A0(_1749_),
    .A1(_1723_),
    .S(net195),
    .X(_3029_));
 sky130_fd_sc_hd__or2_1 _6068_ (.A(net199),
    .B(_3029_),
    .X(_3030_));
 sky130_fd_sc_hd__o21ai_1 _6069_ (.A1(net201),
    .A2(_2970_),
    .B1(_3030_),
    .Y(_3031_));
 sky130_fd_sc_hd__inv_2 _6070_ (.A(_3031_),
    .Y(_3032_));
 sky130_fd_sc_hd__mux2_1 _6071_ (.A0(_2896_),
    .A1(_3031_),
    .S(net207),
    .X(_3033_));
 sky130_fd_sc_hd__or3_1 _6072_ (.A(net210),
    .B(_2851_),
    .C(_3033_),
    .X(_3034_));
 sky130_fd_sc_hd__mux2_1 _6073_ (.A0(_2902_),
    .A1(_2908_),
    .S(net204),
    .X(_3035_));
 sky130_fd_sc_hd__mux2_1 _6074_ (.A0(_2873_),
    .A1(_2906_),
    .S(net206),
    .X(_3036_));
 sky130_fd_sc_hd__mux2_1 _6075_ (.A0(_3035_),
    .A1(_3036_),
    .S(net210),
    .X(_3037_));
 sky130_fd_sc_hd__a21boi_1 _6076_ (.A1(_2821_),
    .A2(_3037_),
    .B1_N(_3034_),
    .Y(_3038_));
 sky130_fd_sc_hd__o221a_1 _6077_ (.A1(_2864_),
    .A2(_3017_),
    .B1(_3038_),
    .B2(net187),
    .C1(_3028_),
    .X(_3039_));
 sky130_fd_sc_hd__o211a_1 _6078_ (.A1(_2861_),
    .A2(_3019_),
    .B1(_3027_),
    .C1(_3039_),
    .X(_3040_));
 sky130_fd_sc_hd__a211oi_1 _6079_ (.A1(_1751_),
    .A2(net224),
    .B1(_3040_),
    .C1(net477),
    .Y(_0819_));
 sky130_fd_sc_hd__a21o_1 _6080_ (.A1(_3016_),
    .A2(_3018_),
    .B1(_3015_),
    .X(_3041_));
 sky130_fd_sc_hd__xnor2_1 _6081_ (.A(_1731_),
    .B(net360),
    .Y(_3042_));
 sky130_fd_sc_hd__nand2_1 _6082_ (.A(_1733_),
    .B(_3042_),
    .Y(_3043_));
 sky130_fd_sc_hd__nor2_1 _6083_ (.A(_1733_),
    .B(_3042_),
    .Y(_3044_));
 sky130_fd_sc_hd__or2_1 _6084_ (.A(_1733_),
    .B(_3042_),
    .X(_3045_));
 sky130_fd_sc_hd__nand2_1 _6085_ (.A(_3043_),
    .B(_3045_),
    .Y(_3046_));
 sky130_fd_sc_hd__a21oi_1 _6086_ (.A1(_3041_),
    .A2(_3046_),
    .B1(net319),
    .Y(_3047_));
 sky130_fd_sc_hd__o21a_1 _6087_ (.A1(_3041_),
    .A2(_3046_),
    .B1(_3047_),
    .X(_3048_));
 sky130_fd_sc_hd__a221o_1 _6088_ (.A1(_1731_),
    .A2(_2857_),
    .B1(_2863_),
    .B2(_1734_),
    .C1(net364),
    .X(_3049_));
 sky130_fd_sc_hd__a21o_1 _6089_ (.A1(_1735_),
    .A2(_3049_),
    .B1(net225),
    .X(_3050_));
 sky130_fd_sc_hd__mux2_1 _6090_ (.A0(_2918_),
    .A1(_2920_),
    .S(net203),
    .X(_3051_));
 sky130_fd_sc_hd__mux2_1 _6091_ (.A0(_2921_),
    .A1(_2931_),
    .S(net203),
    .X(_3052_));
 sky130_fd_sc_hd__or2_1 _6092_ (.A(net209),
    .B(_3051_),
    .X(_3053_));
 sky130_fd_sc_hd__o211a_1 _6093_ (.A1(net213),
    .A2(_3052_),
    .B1(_3053_),
    .C1(_2821_),
    .X(_3054_));
 sky130_fd_sc_hd__mux4_2 _6094_ (.A0(_1723_),
    .A1(_1733_),
    .A2(_1662_),
    .A3(_1749_),
    .S0(net201),
    .S1(net196),
    .X(_3055_));
 sky130_fd_sc_hd__inv_2 _6095_ (.A(_3055_),
    .Y(_3056_));
 sky130_fd_sc_hd__mux2_1 _6096_ (.A0(_2915_),
    .A1(_3056_),
    .S(net206),
    .X(_3057_));
 sky130_fd_sc_hd__or3_1 _6097_ (.A(net209),
    .B(_2851_),
    .C(_3057_),
    .X(_3058_));
 sky130_fd_sc_hd__nand2_1 _6098_ (.A(net189),
    .B(_3058_),
    .Y(_3059_));
 sky130_fd_sc_hd__mux2_1 _6099_ (.A0(_2926_),
    .A1(_2932_),
    .S(net205),
    .X(_3060_));
 sky130_fd_sc_hd__or2_1 _6100_ (.A(net208),
    .B(_3060_),
    .X(_3061_));
 sky130_fd_sc_hd__a21bo_1 _6101_ (.A1(net205),
    .A2(_2936_),
    .B1_N(_2955_),
    .X(_3062_));
 sky130_fd_sc_hd__o21ai_1 _6102_ (.A1(net212),
    .A2(_3062_),
    .B1(_3061_),
    .Y(_3063_));
 sky130_fd_sc_hd__nor2_1 _6103_ (.A(_2817_),
    .B(_3063_),
    .Y(_3064_));
 sky130_fd_sc_hd__nor2_2 _6104_ (.A(net208),
    .B(_2819_),
    .Y(_3065_));
 sky130_fd_sc_hd__nand2_2 _6105_ (.A(net212),
    .B(_2818_),
    .Y(_3066_));
 sky130_fd_sc_hd__or2_1 _6106_ (.A(net202),
    .B(_2928_),
    .X(_3067_));
 sky130_fd_sc_hd__nor2_1 _6107_ (.A(_2819_),
    .B(_3067_),
    .Y(_3068_));
 sky130_fd_sc_hd__o21a_1 _6108_ (.A1(_3065_),
    .A2(_3068_),
    .B1(_3061_),
    .X(_3069_));
 sky130_fd_sc_hd__o32a_2 _6109_ (.A1(net190),
    .A2(_3064_),
    .A3(_3069_),
    .B1(_3054_),
    .B2(_3059_),
    .X(_3070_));
 sky130_fd_sc_hd__nand2_1 _6110_ (.A(_1734_),
    .B(net225),
    .Y(_3071_));
 sky130_fd_sc_hd__o311a_1 _6111_ (.A1(_3048_),
    .A2(_3050_),
    .A3(_3070_),
    .B1(_3071_),
    .C1(net449),
    .X(_0820_));
 sky130_fd_sc_hd__xnor2_1 _6112_ (.A(_1710_),
    .B(net359),
    .Y(_3072_));
 sky130_fd_sc_hd__nor2_1 _6113_ (.A(_1712_),
    .B(_3072_),
    .Y(_3073_));
 sky130_fd_sc_hd__nand2_1 _6114_ (.A(_1712_),
    .B(_3072_),
    .Y(_3074_));
 sky130_fd_sc_hd__nand2b_1 _6115_ (.A_N(_3073_),
    .B(_3074_),
    .Y(_3075_));
 sky130_fd_sc_hd__a21o_2 _6116_ (.A1(_3041_),
    .A2(_3043_),
    .B1(_3044_),
    .X(_3076_));
 sky130_fd_sc_hd__xnor2_1 _6117_ (.A(_3075_),
    .B(_3076_),
    .Y(_3077_));
 sky130_fd_sc_hd__nor2_1 _6118_ (.A(net319),
    .B(_3077_),
    .Y(_3078_));
 sky130_fd_sc_hd__mux4_1 _6119_ (.A0(_1712_),
    .A1(_1733_),
    .A2(_1749_),
    .A3(_1723_),
    .S0(net195),
    .S1(net199),
    .X(_3079_));
 sky130_fd_sc_hd__mux2_1 _6120_ (.A0(_2971_),
    .A1(_3079_),
    .S(net207),
    .X(_3080_));
 sky130_fd_sc_hd__nand2_1 _6121_ (.A(net212),
    .B(_3080_),
    .Y(_3081_));
 sky130_fd_sc_hd__mux2_1 _6122_ (.A0(_2978_),
    .A1(_2980_),
    .S(net203),
    .X(_3082_));
 sky130_fd_sc_hd__mux2_1 _6123_ (.A0(_2950_),
    .A1(_2981_),
    .S(net205),
    .X(_3083_));
 sky130_fd_sc_hd__mux2_1 _6124_ (.A0(_3082_),
    .A1(_3083_),
    .S(net209),
    .X(_3084_));
 sky130_fd_sc_hd__a2bb2o_1 _6125_ (.A1_N(_2851_),
    .A2_N(_3081_),
    .B1(_3084_),
    .B2(_2821_),
    .X(_3085_));
 sky130_fd_sc_hd__o21a_1 _6126_ (.A1(_1710_),
    .A2(_1712_),
    .B1(net363),
    .X(_3086_));
 sky130_fd_sc_hd__a2bb2o_1 _6127_ (.A1_N(_2864_),
    .A2_N(_3075_),
    .B1(_3085_),
    .B2(net189),
    .X(_3087_));
 sky130_fd_sc_hd__a2111o_1 _6128_ (.A1(_1710_),
    .A2(net361),
    .B1(net223),
    .C1(_3086_),
    .D1(_3087_),
    .X(_3088_));
 sky130_fd_sc_hd__mux2_1 _6129_ (.A0(_2951_),
    .A1(_2953_),
    .S(net203),
    .X(_3089_));
 sky130_fd_sc_hd__or2_1 _6130_ (.A(net208),
    .B(_3089_),
    .X(_3090_));
 sky130_fd_sc_hd__o21a_1 _6131_ (.A1(_1467_),
    .A2(net212),
    .B1(_3090_),
    .X(_3091_));
 sky130_fd_sc_hd__and2_1 _6132_ (.A(_2816_),
    .B(_3091_),
    .X(_3092_));
 sky130_fd_sc_hd__nor2_1 _6133_ (.A(net202),
    .B(_2958_),
    .Y(_3093_));
 sky130_fd_sc_hd__o211a_1 _6134_ (.A1(net212),
    .A2(_3093_),
    .B1(_3090_),
    .C1(_2818_),
    .X(_3094_));
 sky130_fd_sc_hd__o21a_1 _6135_ (.A1(_3092_),
    .A2(_3094_),
    .B1(net185),
    .X(_3095_));
 sky130_fd_sc_hd__a21o_1 _6136_ (.A1(_1710_),
    .A2(net2358),
    .B1(net221),
    .X(_3096_));
 sky130_fd_sc_hd__o311a_1 _6137_ (.A1(_3078_),
    .A2(_3088_),
    .A3(_3095_),
    .B1(_3096_),
    .C1(net448),
    .X(_0821_));
 sky130_fd_sc_hd__a21o_1 _6138_ (.A1(_3074_),
    .A2(_3076_),
    .B1(_3073_),
    .X(_3097_));
 sky130_fd_sc_hd__xnor2_1 _6139_ (.A(_1781_),
    .B(net359),
    .Y(_3098_));
 sky130_fd_sc_hd__nand2_1 _6140_ (.A(_1783_),
    .B(_3098_),
    .Y(_3099_));
 sky130_fd_sc_hd__nor2_1 _6141_ (.A(_1783_),
    .B(_3098_),
    .Y(_3100_));
 sky130_fd_sc_hd__inv_2 _6142_ (.A(_3100_),
    .Y(_3101_));
 sky130_fd_sc_hd__nand2_1 _6143_ (.A(_3099_),
    .B(_3101_),
    .Y(_3102_));
 sky130_fd_sc_hd__xnor2_1 _6144_ (.A(_3097_),
    .B(_3102_),
    .Y(_3103_));
 sky130_fd_sc_hd__mux4_1 _6145_ (.A0(_1733_),
    .A1(_1783_),
    .A2(_1749_),
    .A3(_1712_),
    .S0(net201),
    .S1(net195),
    .X(_3104_));
 sky130_fd_sc_hd__mux2_1 _6146_ (.A0(_3006_),
    .A1(_3104_),
    .S(net207),
    .X(_3105_));
 sky130_fd_sc_hd__nand2_1 _6147_ (.A(net214),
    .B(_3105_),
    .Y(_3106_));
 sky130_fd_sc_hd__o31a_1 _6148_ (.A1(net214),
    .A2(net204),
    .A3(_1852_),
    .B1(_3106_),
    .X(_3107_));
 sky130_fd_sc_hd__mux2_1 _6149_ (.A0(_2831_),
    .A1(_2838_),
    .S(net209),
    .X(_3108_));
 sky130_fd_sc_hd__o2bb2a_1 _6150_ (.A1_N(_2821_),
    .A2_N(_3108_),
    .B1(_3107_),
    .B2(_2851_),
    .X(_3109_));
 sky130_fd_sc_hd__nand2_2 _6151_ (.A(_1467_),
    .B(net208),
    .Y(_3110_));
 sky130_fd_sc_hd__nand2_1 _6152_ (.A(net212),
    .B(_2845_),
    .Y(_3111_));
 sky130_fd_sc_hd__o22a_1 _6153_ (.A1(_2817_),
    .A2(_3110_),
    .B1(_3111_),
    .B2(_2820_),
    .X(_3112_));
 sky130_fd_sc_hd__a221o_1 _6154_ (.A1(_1781_),
    .A2(net361),
    .B1(net358),
    .B2(_1784_),
    .C1(net363),
    .X(_3113_));
 sky130_fd_sc_hd__o21ai_1 _6155_ (.A1(_1781_),
    .A2(_1783_),
    .B1(_3113_),
    .Y(_3114_));
 sky130_fd_sc_hd__o211a_1 _6156_ (.A1(net190),
    .A2(_3112_),
    .B1(_3114_),
    .C1(net221),
    .X(_3115_));
 sky130_fd_sc_hd__o221a_1 _6157_ (.A1(net319),
    .A2(_3103_),
    .B1(_3109_),
    .B2(net185),
    .C1(_3115_),
    .X(_3116_));
 sky130_fd_sc_hd__a211oi_1 _6158_ (.A1(_1784_),
    .A2(net223),
    .B1(_3116_),
    .C1(net475),
    .Y(_0822_));
 sky130_fd_sc_hd__xnor2_1 _6159_ (.A(_1760_),
    .B(net360),
    .Y(_3117_));
 sky130_fd_sc_hd__and2_1 _6160_ (.A(_1762_),
    .B(_3117_),
    .X(_3118_));
 sky130_fd_sc_hd__nand2_1 _6161_ (.A(_1762_),
    .B(_3117_),
    .Y(_3119_));
 sky130_fd_sc_hd__nor2_1 _6162_ (.A(_1762_),
    .B(_3117_),
    .Y(_3120_));
 sky130_fd_sc_hd__nor2_1 _6163_ (.A(_3118_),
    .B(_3120_),
    .Y(_3121_));
 sky130_fd_sc_hd__a21o_1 _6164_ (.A1(_3097_),
    .A2(_3099_),
    .B1(_3100_),
    .X(_3122_));
 sky130_fd_sc_hd__nand2_1 _6165_ (.A(_3121_),
    .B(_3122_),
    .Y(_3123_));
 sky130_fd_sc_hd__or2_1 _6166_ (.A(_3121_),
    .B(_3122_),
    .X(_3124_));
 sky130_fd_sc_hd__a21oi_1 _6167_ (.A1(_3123_),
    .A2(_3124_),
    .B1(net2347),
    .Y(_3125_));
 sky130_fd_sc_hd__mux4_1 _6168_ (.A0(_1712_),
    .A1(_1733_),
    .A2(_1762_),
    .A3(_1783_),
    .S0(net195),
    .S1(net201),
    .X(_3126_));
 sky130_fd_sc_hd__mux2_1 _6169_ (.A0(_3032_),
    .A1(_3126_),
    .S(net207),
    .X(_3127_));
 sky130_fd_sc_hd__nor2_1 _6170_ (.A(net210),
    .B(_3127_),
    .Y(_3128_));
 sky130_fd_sc_hd__a211o_1 _6171_ (.A1(net210),
    .A2(_2897_),
    .B1(_3128_),
    .C1(_2851_),
    .X(_3129_));
 sky130_fd_sc_hd__mux2_1 _6172_ (.A0(_2874_),
    .A1(_2909_),
    .S(net213),
    .X(_3130_));
 sky130_fd_sc_hd__nand2_1 _6173_ (.A(_2821_),
    .B(_3130_),
    .Y(_3131_));
 sky130_fd_sc_hd__a21oi_1 _6174_ (.A1(_3129_),
    .A2(_3131_),
    .B1(net186),
    .Y(_3132_));
 sky130_fd_sc_hd__a221o_1 _6175_ (.A1(_1763_),
    .A2(net363),
    .B1(net361),
    .B2(_1760_),
    .C1(net225),
    .X(_3133_));
 sky130_fd_sc_hd__a211o_1 _6176_ (.A1(net358),
    .A2(_3121_),
    .B1(_3132_),
    .C1(_3133_),
    .X(_3134_));
 sky130_fd_sc_hd__mux2_1 _6177_ (.A0(_1468_),
    .A1(_2881_),
    .S(net212),
    .X(_3135_));
 sky130_fd_sc_hd__o2bb2a_1 _6178_ (.A1_N(_2884_),
    .A2_N(_3065_),
    .B1(_3135_),
    .B2(_2817_),
    .X(_3136_));
 sky130_fd_sc_hd__nor2_1 _6179_ (.A(net189),
    .B(_3136_),
    .Y(_3137_));
 sky130_fd_sc_hd__a21o_1 _6180_ (.A1(_1760_),
    .A2(_1762_),
    .B1(net221),
    .X(_3138_));
 sky130_fd_sc_hd__o311a_1 _6181_ (.A1(_3125_),
    .A2(_3134_),
    .A3(_3137_),
    .B1(_3138_),
    .C1(net449),
    .X(_0823_));
 sky130_fd_sc_hd__a21o_1 _6182_ (.A1(_3119_),
    .A2(_3122_),
    .B1(_3120_),
    .X(_3139_));
 sky130_fd_sc_hd__xnor2_1 _6183_ (.A(_1770_),
    .B(net359),
    .Y(_3140_));
 sky130_fd_sc_hd__nand2_1 _6184_ (.A(_1772_),
    .B(_3140_),
    .Y(_3141_));
 sky130_fd_sc_hd__nor2_1 _6185_ (.A(_1772_),
    .B(_3140_),
    .Y(_3142_));
 sky130_fd_sc_hd__or2_1 _6186_ (.A(_1772_),
    .B(_3140_),
    .X(_3143_));
 sky130_fd_sc_hd__nand2_1 _6187_ (.A(_3141_),
    .B(_3143_),
    .Y(_3144_));
 sky130_fd_sc_hd__and2_1 _6188_ (.A(_3139_),
    .B(_3144_),
    .X(_3145_));
 sky130_fd_sc_hd__nor2_1 _6189_ (.A(_3139_),
    .B(_3144_),
    .Y(_3146_));
 sky130_fd_sc_hd__mux4_1 _6190_ (.A0(_1772_),
    .A1(_1783_),
    .A2(_1762_),
    .A3(_1712_),
    .S0(net198),
    .S1(net193),
    .X(_3147_));
 sky130_fd_sc_hd__mux2_1 _6191_ (.A0(_3055_),
    .A1(_3147_),
    .S(net206),
    .X(_3148_));
 sky130_fd_sc_hd__mux2_1 _6192_ (.A0(_2916_),
    .A1(_3148_),
    .S(net213),
    .X(_3149_));
 sky130_fd_sc_hd__nand2_1 _6193_ (.A(_2850_),
    .B(_3149_),
    .Y(_3150_));
 sky130_fd_sc_hd__mux2_1 _6194_ (.A0(_2922_),
    .A1(_2933_),
    .S(net209),
    .X(_3151_));
 sky130_fd_sc_hd__nand2_1 _6195_ (.A(_2821_),
    .B(_3151_),
    .Y(_3152_));
 sky130_fd_sc_hd__a21o_1 _6196_ (.A1(_3150_),
    .A2(_3152_),
    .B1(net186),
    .X(_3153_));
 sky130_fd_sc_hd__a221o_1 _6197_ (.A1(_1770_),
    .A2(net361),
    .B1(net358),
    .B2(_1773_),
    .C1(net363),
    .X(_3154_));
 sky130_fd_sc_hd__o21ai_1 _6198_ (.A1(_1770_),
    .A2(_1772_),
    .B1(_3154_),
    .Y(_3155_));
 sky130_fd_sc_hd__o21a_1 _6199_ (.A1(net208),
    .A2(_2937_),
    .B1(_3110_),
    .X(_3156_));
 sky130_fd_sc_hd__o22a_1 _6200_ (.A1(_2930_),
    .A2(_3066_),
    .B1(_3156_),
    .B2(_2817_),
    .X(_3157_));
 sky130_fd_sc_hd__o211a_1 _6201_ (.A1(net190),
    .A2(_3157_),
    .B1(_3155_),
    .C1(net221),
    .X(_3158_));
 sky130_fd_sc_hd__o311a_1 _6202_ (.A1(net319),
    .A2(_3145_),
    .A3(_3146_),
    .B1(_3153_),
    .C1(_3158_),
    .X(_3159_));
 sky130_fd_sc_hd__a211oi_1 _6203_ (.A1(_1773_),
    .A2(net223),
    .B1(_3159_),
    .C1(net477),
    .Y(_0824_));
 sky130_fd_sc_hd__xnor2_1 _6204_ (.A(_1791_),
    .B(net359),
    .Y(_3160_));
 sky130_fd_sc_hd__and2_1 _6205_ (.A(_1793_),
    .B(_3160_),
    .X(_3161_));
 sky130_fd_sc_hd__nand2_1 _6206_ (.A(_1793_),
    .B(_3160_),
    .Y(_3162_));
 sky130_fd_sc_hd__nor2_1 _6207_ (.A(_1793_),
    .B(_3160_),
    .Y(_3163_));
 sky130_fd_sc_hd__nor2_1 _6208_ (.A(_3161_),
    .B(_3163_),
    .Y(_3164_));
 sky130_fd_sc_hd__a21o_1 _6209_ (.A1(_3139_),
    .A2(_3141_),
    .B1(_3142_),
    .X(_3165_));
 sky130_fd_sc_hd__nand2_1 _6210_ (.A(_3164_),
    .B(_3165_),
    .Y(_3166_));
 sky130_fd_sc_hd__or2_1 _6211_ (.A(_3164_),
    .B(_3165_),
    .X(_3167_));
 sky130_fd_sc_hd__a21oi_1 _6212_ (.A1(_3166_),
    .A2(_3167_),
    .B1(net319),
    .Y(_3168_));
 sky130_fd_sc_hd__mux4_1 _6213_ (.A0(_1762_),
    .A1(_1783_),
    .A2(_1793_),
    .A3(_1772_),
    .S0(net193),
    .S1(net200),
    .X(_3169_));
 sky130_fd_sc_hd__mux2_1 _6214_ (.A0(_3079_),
    .A1(_3169_),
    .S(net207),
    .X(_3170_));
 sky130_fd_sc_hd__nor2_1 _6215_ (.A(net210),
    .B(_3170_),
    .Y(_3171_));
 sky130_fd_sc_hd__a211o_1 _6216_ (.A1(net210),
    .A2(_2972_),
    .B1(_3171_),
    .C1(_2851_),
    .X(_3172_));
 sky130_fd_sc_hd__mux2_1 _6217_ (.A0(_2952_),
    .A1(_2982_),
    .S(net213),
    .X(_3173_));
 sky130_fd_sc_hd__a21bo_1 _6218_ (.A1(_2821_),
    .A2(_3173_),
    .B1_N(_3172_),
    .X(_3174_));
 sky130_fd_sc_hd__a221o_1 _6219_ (.A1(_1794_),
    .A2(net364),
    .B1(net362),
    .B2(_1791_),
    .C1(net225),
    .X(_3175_));
 sky130_fd_sc_hd__a22o_1 _6220_ (.A1(net358),
    .A2(_3164_),
    .B1(_3174_),
    .B2(net190),
    .X(_3176_));
 sky130_fd_sc_hd__a21bo_1 _6221_ (.A1(net212),
    .A2(_2956_),
    .B1_N(_3110_),
    .X(_3177_));
 sky130_fd_sc_hd__a22o_1 _6222_ (.A1(_2960_),
    .A2(_3065_),
    .B1(_3177_),
    .B2(_2816_),
    .X(_3178_));
 sky130_fd_sc_hd__a211o_1 _6223_ (.A1(net185),
    .A2(_3178_),
    .B1(_3176_),
    .C1(_3175_),
    .X(_3179_));
 sky130_fd_sc_hd__a21o_1 _6224_ (.A1(_1791_),
    .A2(net2362),
    .B1(net221),
    .X(_3180_));
 sky130_fd_sc_hd__o211a_1 _6225_ (.A1(_3168_),
    .A2(_3179_),
    .B1(_3180_),
    .C1(net448),
    .X(_0825_));
 sky130_fd_sc_hd__a21o_2 _6226_ (.A1(_3162_),
    .A2(_3165_),
    .B1(_3163_),
    .X(_3181_));
 sky130_fd_sc_hd__xnor2_1 _6227_ (.A(_1825_),
    .B(net360),
    .Y(_3182_));
 sky130_fd_sc_hd__nand2_1 _6228_ (.A(_1828_),
    .B(_3182_),
    .Y(_3183_));
 sky130_fd_sc_hd__nor2_1 _6229_ (.A(_1828_),
    .B(_3182_),
    .Y(_3184_));
 sky130_fd_sc_hd__or2_1 _6230_ (.A(_1828_),
    .B(_3182_),
    .X(_3185_));
 sky130_fd_sc_hd__nand2_1 _6231_ (.A(_3183_),
    .B(_3185_),
    .Y(_3186_));
 sky130_fd_sc_hd__o21ai_1 _6232_ (.A1(_3181_),
    .A2(_3186_),
    .B1(_2862_),
    .Y(_3187_));
 sky130_fd_sc_hd__a21oi_1 _6233_ (.A1(_3181_),
    .A2(_3186_),
    .B1(_3187_),
    .Y(_3188_));
 sky130_fd_sc_hd__mux4_1 _6234_ (.A0(_1772_),
    .A1(_1828_),
    .A2(_1762_),
    .A3(_1793_),
    .S0(net201),
    .S1(net195),
    .X(_3189_));
 sky130_fd_sc_hd__mux2_1 _6235_ (.A0(_3104_),
    .A1(_3189_),
    .S(net207),
    .X(_3190_));
 sky130_fd_sc_hd__nand2_1 _6236_ (.A(net211),
    .B(_3008_),
    .Y(_3191_));
 sky130_fd_sc_hd__o211a_1 _6237_ (.A1(net211),
    .A2(_3190_),
    .B1(_3191_),
    .C1(_2850_),
    .X(_3192_));
 sky130_fd_sc_hd__or2_1 _6238_ (.A(net208),
    .B(_3001_),
    .X(_3193_));
 sky130_fd_sc_hd__o211a_1 _6239_ (.A1(net214),
    .A2(_2995_),
    .B1(_3193_),
    .C1(_2821_),
    .X(_3194_));
 sky130_fd_sc_hd__o21a_1 _6240_ (.A1(_3192_),
    .A2(_3194_),
    .B1(net191),
    .X(_3195_));
 sky130_fd_sc_hd__a2bb2o_1 _6241_ (.A1_N(_2864_),
    .A2_N(_1829_),
    .B1(_1825_),
    .B2(net362),
    .X(_3196_));
 sky130_fd_sc_hd__o21ba_1 _6242_ (.A1(net364),
    .A2(_3196_),
    .B1_N(_1830_),
    .X(_3197_));
 sky130_fd_sc_hd__o21ai_1 _6243_ (.A1(net208),
    .A2(_2997_),
    .B1(_3110_),
    .Y(_3198_));
 sky130_fd_sc_hd__a22o_2 _6244_ (.A1(_2996_),
    .A2(_3065_),
    .B1(_3198_),
    .B2(_2816_),
    .X(_3199_));
 sky130_fd_sc_hd__a2111o_1 _6245_ (.A1(net188),
    .A2(_3199_),
    .B1(_3197_),
    .C1(_3195_),
    .D1(net224),
    .X(_3200_));
 sky130_fd_sc_hd__o221a_1 _6246_ (.A1(_1829_),
    .A2(net222),
    .B1(_3188_),
    .B2(_3200_),
    .C1(net461),
    .X(_0826_));
 sky130_fd_sc_hd__xnor2_1 _6247_ (.A(_1803_),
    .B(net360),
    .Y(_3201_));
 sky130_fd_sc_hd__and2_1 _6248_ (.A(_1806_),
    .B(_3201_),
    .X(_3202_));
 sky130_fd_sc_hd__nand2_1 _6249_ (.A(_1806_),
    .B(_3201_),
    .Y(_3203_));
 sky130_fd_sc_hd__nor2_1 _6250_ (.A(_1806_),
    .B(_3201_),
    .Y(_3204_));
 sky130_fd_sc_hd__nor2_1 _6251_ (.A(_3202_),
    .B(_3204_),
    .Y(_3205_));
 sky130_fd_sc_hd__a21o_1 _6252_ (.A1(_3181_),
    .A2(_3183_),
    .B1(_3184_),
    .X(_3206_));
 sky130_fd_sc_hd__xnor2_1 _6253_ (.A(_3205_),
    .B(_3206_),
    .Y(_3207_));
 sky130_fd_sc_hd__mux4_1 _6254_ (.A0(_1793_),
    .A1(_1806_),
    .A2(_1772_),
    .A3(_1828_),
    .S0(net201),
    .S1(net195),
    .X(_3208_));
 sky130_fd_sc_hd__mux2_1 _6255_ (.A0(_3126_),
    .A1(_3208_),
    .S(net207),
    .X(_3209_));
 sky130_fd_sc_hd__nor2_1 _6256_ (.A(net210),
    .B(_3209_),
    .Y(_3210_));
 sky130_fd_sc_hd__a211o_1 _6257_ (.A1(net210),
    .A2(_3033_),
    .B1(_3210_),
    .C1(_2851_),
    .X(_3211_));
 sky130_fd_sc_hd__mux2_1 _6258_ (.A0(_3020_),
    .A1(_3036_),
    .S(net214),
    .X(_3212_));
 sky130_fd_sc_hd__a21bo_1 _6259_ (.A1(_2821_),
    .A2(_3212_),
    .B1_N(_3211_),
    .X(_3213_));
 sky130_fd_sc_hd__o21a_1 _6260_ (.A1(_1803_),
    .A2(_1806_),
    .B1(net364),
    .X(_3214_));
 sky130_fd_sc_hd__a22o_1 _6261_ (.A1(_2863_),
    .A2(_3205_),
    .B1(_3213_),
    .B2(net191),
    .X(_3215_));
 sky130_fd_sc_hd__a2111o_1 _6262_ (.A1(_1803_),
    .A2(net362),
    .B1(net225),
    .C1(_3214_),
    .D1(_3215_),
    .X(_3216_));
 sky130_fd_sc_hd__o21a_1 _6263_ (.A1(net208),
    .A2(_3022_),
    .B1(_3110_),
    .X(_3217_));
 sky130_fd_sc_hd__o22ai_4 _6264_ (.A1(_3025_),
    .A2(_3066_),
    .B1(_3217_),
    .B2(_2817_),
    .Y(_3218_));
 sky130_fd_sc_hd__a22o_1 _6265_ (.A1(_2862_),
    .A2(_3207_),
    .B1(_3218_),
    .B2(net188),
    .X(_3219_));
 sky130_fd_sc_hd__a21o_1 _6266_ (.A1(_1803_),
    .A2(_1806_),
    .B1(net222),
    .X(_3220_));
 sky130_fd_sc_hd__o211a_1 _6267_ (.A1(_3216_),
    .A2(_3219_),
    .B1(_3220_),
    .C1(net461),
    .X(_0827_));
 sky130_fd_sc_hd__a21o_1 _6268_ (.A1(_3203_),
    .A2(_3206_),
    .B1(_3204_),
    .X(_3221_));
 sky130_fd_sc_hd__xnor2_1 _6269_ (.A(_1813_),
    .B(net360),
    .Y(_3222_));
 sky130_fd_sc_hd__nand2_1 _6270_ (.A(_1815_),
    .B(_3222_),
    .Y(_3223_));
 sky130_fd_sc_hd__nor2_1 _6271_ (.A(_1815_),
    .B(_3222_),
    .Y(_3224_));
 sky130_fd_sc_hd__or2_1 _6272_ (.A(_1815_),
    .B(_3222_),
    .X(_3225_));
 sky130_fd_sc_hd__nand2_1 _6273_ (.A(_3223_),
    .B(_3225_),
    .Y(_3226_));
 sky130_fd_sc_hd__or2_1 _6274_ (.A(_3221_),
    .B(_3226_),
    .X(_3227_));
 sky130_fd_sc_hd__nand2_1 _6275_ (.A(_3221_),
    .B(_3226_),
    .Y(_3228_));
 sky130_fd_sc_hd__mux4_1 _6276_ (.A0(_1815_),
    .A1(_1828_),
    .A2(_1806_),
    .A3(_1793_),
    .S0(net198),
    .S1(net193),
    .X(_3229_));
 sky130_fd_sc_hd__or2_1 _6277_ (.A(net205),
    .B(_3147_),
    .X(_3230_));
 sky130_fd_sc_hd__o21ai_1 _6278_ (.A1(net203),
    .A2(_3229_),
    .B1(_3230_),
    .Y(_3231_));
 sky130_fd_sc_hd__and2_1 _6279_ (.A(net213),
    .B(_3231_),
    .X(_3232_));
 sky130_fd_sc_hd__a211o_1 _6280_ (.A1(net209),
    .A2(_3057_),
    .B1(_3232_),
    .C1(_2851_),
    .X(_3233_));
 sky130_fd_sc_hd__mux2_1 _6281_ (.A0(_3052_),
    .A1(_3060_),
    .S(net209),
    .X(_3234_));
 sky130_fd_sc_hd__a21bo_2 _6282_ (.A1(_2821_),
    .A2(_3234_),
    .B1_N(_3233_),
    .X(_3235_));
 sky130_fd_sc_hd__a2bb2o_1 _6283_ (.A1_N(_2864_),
    .A2_N(_1816_),
    .B1(_1813_),
    .B2(net362),
    .X(_3236_));
 sky130_fd_sc_hd__o21ba_1 _6284_ (.A1(net364),
    .A2(_3236_),
    .B1_N(_1817_),
    .X(_3237_));
 sky130_fd_sc_hd__a21bo_1 _6285_ (.A1(net212),
    .A2(_3062_),
    .B1_N(_3110_),
    .X(_3238_));
 sky130_fd_sc_hd__a22o_2 _6286_ (.A1(net212),
    .A2(_3068_),
    .B1(_3238_),
    .B2(_2816_),
    .X(_3239_));
 sky130_fd_sc_hd__a211o_1 _6287_ (.A1(net191),
    .A2(_3235_),
    .B1(_3237_),
    .C1(net224),
    .X(_3240_));
 sky130_fd_sc_hd__a32o_1 _6288_ (.A1(_2862_),
    .A2(_3227_),
    .A3(_3228_),
    .B1(_3239_),
    .B2(net188),
    .X(_3241_));
 sky130_fd_sc_hd__o221a_1 _6289_ (.A1(_1816_),
    .A2(net222),
    .B1(_3240_),
    .B2(_3241_),
    .C1(net459),
    .X(_0828_));
 sky130_fd_sc_hd__xnor2_1 _6290_ (.A(_1837_),
    .B(net360),
    .Y(_3242_));
 sky130_fd_sc_hd__and2_1 _6291_ (.A(_1839_),
    .B(_3242_),
    .X(_3243_));
 sky130_fd_sc_hd__nand2_1 _6292_ (.A(_1839_),
    .B(_3242_),
    .Y(_3244_));
 sky130_fd_sc_hd__nor2_1 _6293_ (.A(_1839_),
    .B(_3242_),
    .Y(_3245_));
 sky130_fd_sc_hd__nor2_1 _6294_ (.A(_3243_),
    .B(_3245_),
    .Y(_3246_));
 sky130_fd_sc_hd__a21o_1 _6295_ (.A1(_3221_),
    .A2(_3223_),
    .B1(_3224_),
    .X(_3247_));
 sky130_fd_sc_hd__nand2_1 _6296_ (.A(_3246_),
    .B(_3247_),
    .Y(_3248_));
 sky130_fd_sc_hd__or2_1 _6297_ (.A(_3246_),
    .B(_3247_),
    .X(_3249_));
 sky130_fd_sc_hd__a21oi_1 _6298_ (.A1(_3248_),
    .A2(_3249_),
    .B1(net2347),
    .Y(_3250_));
 sky130_fd_sc_hd__mux4_1 _6299_ (.A0(_1806_),
    .A1(_1828_),
    .A2(_1839_),
    .A3(_1815_),
    .S0(net193),
    .S1(net200),
    .X(_3251_));
 sky130_fd_sc_hd__mux2_1 _6300_ (.A0(_3169_),
    .A1(_3251_),
    .S(net206),
    .X(_3252_));
 sky130_fd_sc_hd__mux2_2 _6301_ (.A0(_3080_),
    .A1(_3252_),
    .S(net213),
    .X(_3253_));
 sky130_fd_sc_hd__a221o_1 _6302_ (.A1(_1840_),
    .A2(net364),
    .B1(net362),
    .B2(_1837_),
    .C1(net224),
    .X(_3254_));
 sky130_fd_sc_hd__a221o_1 _6303_ (.A1(_2863_),
    .A2(_3246_),
    .B1(_3253_),
    .B2(_2852_),
    .C1(_3254_),
    .X(_3255_));
 sky130_fd_sc_hd__o21a_4 _6304_ (.A1(_1467_),
    .A2(net189),
    .B1(_2816_),
    .X(_3256_));
 sky130_fd_sc_hd__o21ai_4 _6305_ (.A1(_1467_),
    .A2(net189),
    .B1(_2816_),
    .Y(_3257_));
 sky130_fd_sc_hd__nand2_1 _6306_ (.A(net212),
    .B(_3093_),
    .Y(_3258_));
 sky130_fd_sc_hd__a21oi_1 _6307_ (.A1(net185),
    .A2(_3258_),
    .B1(_2819_),
    .Y(_3259_));
 sky130_fd_sc_hd__mux2_1 _6308_ (.A0(_3083_),
    .A1(_3089_),
    .S(net208),
    .X(_3260_));
 sky130_fd_sc_hd__o22a_2 _6309_ (.A1(_3256_),
    .A2(_3259_),
    .B1(_3260_),
    .B2(net186),
    .X(_3261_));
 sky130_fd_sc_hd__a21oi_1 _6310_ (.A1(_1841_),
    .A2(net224),
    .B1(net477),
    .Y(_3262_));
 sky130_fd_sc_hd__o31a_1 _6311_ (.A1(_3250_),
    .A2(_3255_),
    .A3(_3261_),
    .B1(_3262_),
    .X(_0829_));
 sky130_fd_sc_hd__a21o_1 _6312_ (.A1(_3244_),
    .A2(_3247_),
    .B1(_3245_),
    .X(_3263_));
 sky130_fd_sc_hd__xnor2_1 _6313_ (.A(_1541_),
    .B(_2859_),
    .Y(_3264_));
 sky130_fd_sc_hd__nand2_1 _6314_ (.A(_1544_),
    .B(_3264_),
    .Y(_3265_));
 sky130_fd_sc_hd__nor2_1 _6315_ (.A(_1544_),
    .B(_3264_),
    .Y(_3266_));
 sky130_fd_sc_hd__or2_1 _6316_ (.A(_1544_),
    .B(_3264_),
    .X(_3267_));
 sky130_fd_sc_hd__nand2_1 _6317_ (.A(_3265_),
    .B(_3267_),
    .Y(_3268_));
 sky130_fd_sc_hd__and2_1 _6318_ (.A(_3263_),
    .B(_3268_),
    .X(_3269_));
 sky130_fd_sc_hd__nor2_1 _6319_ (.A(_3263_),
    .B(_3268_),
    .Y(_3270_));
 sky130_fd_sc_hd__nand2_1 _6320_ (.A(net210),
    .B(_3105_),
    .Y(_3271_));
 sky130_fd_sc_hd__mux4_1 _6321_ (.A0(_1544_),
    .A1(_1815_),
    .A2(_1839_),
    .A3(_1806_),
    .S0(net198),
    .S1(net195),
    .X(_3272_));
 sky130_fd_sc_hd__mux2_1 _6322_ (.A0(_3189_),
    .A1(_3272_),
    .S(net206),
    .X(_3273_));
 sky130_fd_sc_hd__a21oi_1 _6323_ (.A1(net214),
    .A2(_3273_),
    .B1(net187),
    .Y(_3274_));
 sky130_fd_sc_hd__a221o_1 _6324_ (.A1(net187),
    .A2(_2849_),
    .B1(_3271_),
    .B2(_3274_),
    .C1(_2851_),
    .X(_3275_));
 sky130_fd_sc_hd__nor2_2 _6325_ (.A(net185),
    .B(_2819_),
    .Y(_3276_));
 sky130_fd_sc_hd__a221o_1 _6326_ (.A1(_1542_),
    .A2(net362),
    .B1(net358),
    .B2(_1545_),
    .C1(net364),
    .X(_3277_));
 sky130_fd_sc_hd__o21a_1 _6327_ (.A1(_1542_),
    .A2(_1544_),
    .B1(_3277_),
    .X(_3278_));
 sky130_fd_sc_hd__o21a_1 _6328_ (.A1(net187),
    .A2(_2846_),
    .B1(_3256_),
    .X(_3279_));
 sky130_fd_sc_hd__a2111oi_1 _6329_ (.A1(_2846_),
    .A2(_3276_),
    .B1(_3278_),
    .C1(_3279_),
    .D1(net224),
    .Y(_3280_));
 sky130_fd_sc_hd__o311a_1 _6330_ (.A1(net319),
    .A2(_3269_),
    .A3(_3270_),
    .B1(_3275_),
    .C1(_3280_),
    .X(_3281_));
 sky130_fd_sc_hd__a211oi_1 _6331_ (.A1(_1545_),
    .A2(net224),
    .B1(_3281_),
    .C1(net477),
    .Y(_0830_));
 sky130_fd_sc_hd__xnor2_2 _6332_ (.A(_1518_),
    .B(net360),
    .Y(_3282_));
 sky130_fd_sc_hd__nand2_1 _6333_ (.A(_1521_),
    .B(_3282_),
    .Y(_3283_));
 sky130_fd_sc_hd__nor2_1 _6334_ (.A(_1521_),
    .B(_3282_),
    .Y(_3284_));
 sky130_fd_sc_hd__xnor2_1 _6335_ (.A(_1520_),
    .B(_3282_),
    .Y(_3285_));
 sky130_fd_sc_hd__a21o_1 _6336_ (.A1(_3263_),
    .A2(_3265_),
    .B1(_3266_),
    .X(_3286_));
 sky130_fd_sc_hd__xnor2_1 _6337_ (.A(_3285_),
    .B(_3286_),
    .Y(_3287_));
 sky130_fd_sc_hd__mux4_1 _6338_ (.A0(_1521_),
    .A1(_1544_),
    .A2(_1839_),
    .A3(_1815_),
    .S0(net195),
    .S1(net198),
    .X(_3288_));
 sky130_fd_sc_hd__mux2_1 _6339_ (.A0(_3208_),
    .A1(_3288_),
    .S(net206),
    .X(_3289_));
 sky130_fd_sc_hd__mux2_1 _6340_ (.A0(_3127_),
    .A1(_3289_),
    .S(net214),
    .X(_3290_));
 sky130_fd_sc_hd__nand2_1 _6341_ (.A(net187),
    .B(_2898_),
    .Y(_3291_));
 sky130_fd_sc_hd__o211a_1 _6342_ (.A1(net187),
    .A2(_3290_),
    .B1(_3291_),
    .C1(_2850_),
    .X(_3292_));
 sky130_fd_sc_hd__a221o_1 _6343_ (.A1(_1522_),
    .A2(net364),
    .B1(net362),
    .B2(_1518_),
    .C1(net224),
    .X(_3293_));
 sky130_fd_sc_hd__a221o_1 _6344_ (.A1(_2885_),
    .A2(_3276_),
    .B1(_3285_),
    .B2(net358),
    .C1(_3293_),
    .X(_3294_));
 sky130_fd_sc_hd__or2_1 _6345_ (.A(net188),
    .B(_2882_),
    .X(_3295_));
 sky130_fd_sc_hd__a22o_1 _6346_ (.A1(_2862_),
    .A2(_3287_),
    .B1(_3295_),
    .B2(_3256_),
    .X(_3296_));
 sky130_fd_sc_hd__nand2_1 _6347_ (.A(_1523_),
    .B(net224),
    .Y(_3297_));
 sky130_fd_sc_hd__o311a_1 _6348_ (.A1(_3292_),
    .A2(_3294_),
    .A3(_3296_),
    .B1(_3297_),
    .C1(net453),
    .X(_0831_));
 sky130_fd_sc_hd__a21o_1 _6349_ (.A1(_3283_),
    .A2(_3286_),
    .B1(_3284_),
    .X(_3298_));
 sky130_fd_sc_hd__xnor2_1 _6350_ (.A(_1553_),
    .B(net360),
    .Y(_3299_));
 sky130_fd_sc_hd__nand2_1 _6351_ (.A(_1555_),
    .B(_3299_),
    .Y(_3300_));
 sky130_fd_sc_hd__nor2_1 _6352_ (.A(_1555_),
    .B(_3299_),
    .Y(_3301_));
 sky130_fd_sc_hd__or2_1 _6353_ (.A(_1555_),
    .B(_3299_),
    .X(_3302_));
 sky130_fd_sc_hd__nand2_1 _6354_ (.A(_3300_),
    .B(_3302_),
    .Y(_3303_));
 sky130_fd_sc_hd__or2_1 _6355_ (.A(_3298_),
    .B(_3303_),
    .X(_3304_));
 sky130_fd_sc_hd__nand2_1 _6356_ (.A(_3298_),
    .B(_3303_),
    .Y(_3305_));
 sky130_fd_sc_hd__a21oi_1 _6357_ (.A1(_1468_),
    .A2(net186),
    .B1(_2938_),
    .Y(_3306_));
 sky130_fd_sc_hd__a221o_1 _6358_ (.A1(_1553_),
    .A2(net362),
    .B1(_2863_),
    .B2(_1556_),
    .C1(_2856_),
    .X(_3307_));
 sky130_fd_sc_hd__a32o_1 _6359_ (.A1(net214),
    .A2(_2850_),
    .A3(_2916_),
    .B1(_2816_),
    .B2(_1467_),
    .X(_3308_));
 sky130_fd_sc_hd__a221o_1 _6360_ (.A1(_1557_),
    .A2(_3307_),
    .B1(_3308_),
    .B2(net188),
    .C1(net224),
    .X(_3309_));
 sky130_fd_sc_hd__mux4_1 _6361_ (.A0(_1544_),
    .A1(_1839_),
    .A2(_1555_),
    .A3(_1521_),
    .S0(net193),
    .S1(net200),
    .X(_3310_));
 sky130_fd_sc_hd__mux2_1 _6362_ (.A0(_3229_),
    .A1(_3310_),
    .S(net205),
    .X(_3311_));
 sky130_fd_sc_hd__mux2_1 _6363_ (.A0(_3148_),
    .A1(_3311_),
    .S(net213),
    .X(_3312_));
 sky130_fd_sc_hd__a21bo_1 _6364_ (.A1(_2850_),
    .A2(_3312_),
    .B1_N(_2935_),
    .X(_3313_));
 sky130_fd_sc_hd__a32o_1 _6365_ (.A1(_2862_),
    .A2(_3304_),
    .A3(_3305_),
    .B1(_3313_),
    .B2(net191),
    .X(_3314_));
 sky130_fd_sc_hd__a21oi_1 _6366_ (.A1(_1556_),
    .A2(net225),
    .B1(net477),
    .Y(_3315_));
 sky130_fd_sc_hd__o31a_1 _6367_ (.A1(_3306_),
    .A2(_3309_),
    .A3(_3314_),
    .B1(_3315_),
    .X(_0832_));
 sky130_fd_sc_hd__xnor2_1 _6368_ (.A(_1529_),
    .B(net360),
    .Y(_3316_));
 sky130_fd_sc_hd__and2_1 _6369_ (.A(_1531_),
    .B(_3316_),
    .X(_3317_));
 sky130_fd_sc_hd__nand2_1 _6370_ (.A(_1531_),
    .B(_3316_),
    .Y(_3318_));
 sky130_fd_sc_hd__nor2_1 _6371_ (.A(_1531_),
    .B(_3316_),
    .Y(_3319_));
 sky130_fd_sc_hd__nor2_1 _6372_ (.A(_3317_),
    .B(_3319_),
    .Y(_3320_));
 sky130_fd_sc_hd__a21o_1 _6373_ (.A1(_3298_),
    .A2(_3300_),
    .B1(_3301_),
    .X(_3321_));
 sky130_fd_sc_hd__xnor2_1 _6374_ (.A(_3320_),
    .B(_3321_),
    .Y(_3322_));
 sky130_fd_sc_hd__mux4_1 _6375_ (.A0(_1521_),
    .A1(_1531_),
    .A2(_1544_),
    .A3(_1555_),
    .S0(net200),
    .S1(net194),
    .X(_3323_));
 sky130_fd_sc_hd__mux2_1 _6376_ (.A0(_3251_),
    .A1(_3323_),
    .S(net206),
    .X(_3324_));
 sky130_fd_sc_hd__mux2_1 _6377_ (.A0(_3170_),
    .A1(_3324_),
    .S(net214),
    .X(_3325_));
 sky130_fd_sc_hd__nand2_1 _6378_ (.A(net187),
    .B(_2973_),
    .Y(_3326_));
 sky130_fd_sc_hd__o211a_1 _6379_ (.A1(net187),
    .A2(_3325_),
    .B1(_3326_),
    .C1(_2850_),
    .X(_3327_));
 sky130_fd_sc_hd__a221o_1 _6380_ (.A1(_1532_),
    .A2(net364),
    .B1(net362),
    .B2(_1529_),
    .C1(net224),
    .X(_3328_));
 sky130_fd_sc_hd__a221o_1 _6381_ (.A1(_2961_),
    .A2(_3276_),
    .B1(_3320_),
    .B2(_2863_),
    .C1(_3328_),
    .X(_3329_));
 sky130_fd_sc_hd__or2_1 _6382_ (.A(net187),
    .B(_2957_),
    .X(_3330_));
 sky130_fd_sc_hd__a221o_1 _6383_ (.A1(_2862_),
    .A2(_3322_),
    .B1(_3330_),
    .B2(_3256_),
    .C1(_3329_),
    .X(_3331_));
 sky130_fd_sc_hd__a21o_1 _6384_ (.A1(_1529_),
    .A2(net2367),
    .B1(net222),
    .X(_3332_));
 sky130_fd_sc_hd__o211a_1 _6385_ (.A1(_3327_),
    .A2(_3331_),
    .B1(_3332_),
    .C1(net453),
    .X(_0833_));
 sky130_fd_sc_hd__a21o_1 _6386_ (.A1(_3318_),
    .A2(_3321_),
    .B1(_3319_),
    .X(_3333_));
 sky130_fd_sc_hd__xnor2_1 _6387_ (.A(_1588_),
    .B(net359),
    .Y(_3334_));
 sky130_fd_sc_hd__and2_1 _6388_ (.A(_1590_),
    .B(_3334_),
    .X(_3335_));
 sky130_fd_sc_hd__nand2_1 _6389_ (.A(_1590_),
    .B(_3334_),
    .Y(_3336_));
 sky130_fd_sc_hd__nor2_1 _6390_ (.A(_1590_),
    .B(_3334_),
    .Y(_3337_));
 sky130_fd_sc_hd__nor2_1 _6391_ (.A(_3335_),
    .B(_3337_),
    .Y(_3338_));
 sky130_fd_sc_hd__xnor2_1 _6392_ (.A(_3333_),
    .B(_3338_),
    .Y(_3339_));
 sky130_fd_sc_hd__mux4_1 _6393_ (.A0(_1590_),
    .A1(_1555_),
    .A2(_1531_),
    .A3(_1521_),
    .S0(net198),
    .S1(net194),
    .X(_3340_));
 sky130_fd_sc_hd__mux2_1 _6394_ (.A0(_3272_),
    .A1(_3340_),
    .S(net206),
    .X(_3341_));
 sky130_fd_sc_hd__o21a_1 _6395_ (.A1(net212),
    .A2(_2996_),
    .B1(_3276_),
    .X(_3342_));
 sky130_fd_sc_hd__o22a_1 _6396_ (.A1(net185),
    .A2(_2999_),
    .B1(_3256_),
    .B2(_3342_),
    .X(_3343_));
 sky130_fd_sc_hd__a221o_1 _6397_ (.A1(_1588_),
    .A2(net361),
    .B1(net358),
    .B2(_1591_),
    .C1(net363),
    .X(_3344_));
 sky130_fd_sc_hd__o21a_1 _6398_ (.A1(_1588_),
    .A2(_1590_),
    .B1(_3344_),
    .X(_3345_));
 sky130_fd_sc_hd__o2bb2a_1 _6399_ (.A1_N(net187),
    .A2_N(_3009_),
    .B1(_3190_),
    .B2(net214),
    .X(_3346_));
 sky130_fd_sc_hd__o311a_1 _6400_ (.A1(net210),
    .A2(net187),
    .A3(_3341_),
    .B1(_3346_),
    .C1(_2850_),
    .X(_3347_));
 sky130_fd_sc_hd__or4_1 _6401_ (.A(net223),
    .B(_3343_),
    .C(_3345_),
    .D(_3347_),
    .X(_3348_));
 sky130_fd_sc_hd__a21oi_1 _6402_ (.A1(_2862_),
    .A2(_3339_),
    .B1(_3348_),
    .Y(_3349_));
 sky130_fd_sc_hd__a211oi_1 _6403_ (.A1(net2316),
    .A2(net223),
    .B1(_3349_),
    .C1(net473),
    .Y(_0834_));
 sky130_fd_sc_hd__xnor2_1 _6404_ (.A(_1565_),
    .B(net359),
    .Y(_3350_));
 sky130_fd_sc_hd__and2_1 _6405_ (.A(_1567_),
    .B(_3350_),
    .X(_3351_));
 sky130_fd_sc_hd__nand2_1 _6406_ (.A(_1567_),
    .B(_3350_),
    .Y(_3352_));
 sky130_fd_sc_hd__nor2_1 _6407_ (.A(_1567_),
    .B(_3350_),
    .Y(_3353_));
 sky130_fd_sc_hd__nor2_1 _6408_ (.A(_3351_),
    .B(_3353_),
    .Y(_3354_));
 sky130_fd_sc_hd__a21o_1 _6409_ (.A1(_3333_),
    .A2(_3336_),
    .B1(_3337_),
    .X(_3355_));
 sky130_fd_sc_hd__xnor2_1 _6410_ (.A(_3354_),
    .B(_3355_),
    .Y(_3356_));
 sky130_fd_sc_hd__a21oi_1 _6411_ (.A1(net189),
    .A2(_3023_),
    .B1(_3257_),
    .Y(_3357_));
 sky130_fd_sc_hd__a221o_1 _6412_ (.A1(_1568_),
    .A2(net363),
    .B1(net361),
    .B2(_1565_),
    .C1(net223),
    .X(_3358_));
 sky130_fd_sc_hd__a221o_1 _6413_ (.A1(net189),
    .A2(_3026_),
    .B1(_3354_),
    .B2(net358),
    .C1(_3358_),
    .X(_3359_));
 sky130_fd_sc_hd__mux4_1 _6414_ (.A0(_1531_),
    .A1(_1555_),
    .A2(_1567_),
    .A3(_1590_),
    .S0(net194),
    .S1(net200),
    .X(_3360_));
 sky130_fd_sc_hd__mux2_1 _6415_ (.A0(_3288_),
    .A1(_3360_),
    .S(net206),
    .X(_3361_));
 sky130_fd_sc_hd__mux2_1 _6416_ (.A0(_3209_),
    .A1(_3361_),
    .S(net214),
    .X(_3362_));
 sky130_fd_sc_hd__o2bb2a_1 _6417_ (.A1_N(_2853_),
    .A2_N(_3034_),
    .B1(_3362_),
    .B2(net187),
    .X(_3363_));
 sky130_fd_sc_hd__a21o_1 _6418_ (.A1(_2862_),
    .A2(_3356_),
    .B1(_3363_),
    .X(_3364_));
 sky130_fd_sc_hd__a21o_1 _6419_ (.A1(_1565_),
    .A2(_1567_),
    .B1(net221),
    .X(_3365_));
 sky130_fd_sc_hd__o311a_1 _6420_ (.A1(_3357_),
    .A2(_3359_),
    .A3(_3364_),
    .B1(_3365_),
    .C1(net454),
    .X(_0835_));
 sky130_fd_sc_hd__a21o_1 _6421_ (.A1(_3352_),
    .A2(_3355_),
    .B1(_3353_),
    .X(_3366_));
 sky130_fd_sc_hd__xnor2_1 _6422_ (.A(_1575_),
    .B(net359),
    .Y(_3367_));
 sky130_fd_sc_hd__nand2_1 _6423_ (.A(_1577_),
    .B(_3367_),
    .Y(_3368_));
 sky130_fd_sc_hd__nor2_1 _6424_ (.A(_1577_),
    .B(_3367_),
    .Y(_3369_));
 sky130_fd_sc_hd__or2_1 _6425_ (.A(_1577_),
    .B(_3367_),
    .X(_3370_));
 sky130_fd_sc_hd__nand2_1 _6426_ (.A(_3368_),
    .B(_3370_),
    .Y(_3371_));
 sky130_fd_sc_hd__xnor2_1 _6427_ (.A(_3366_),
    .B(_3371_),
    .Y(_3372_));
 sky130_fd_sc_hd__mux4_1 _6428_ (.A0(_1577_),
    .A1(_1590_),
    .A2(_1567_),
    .A3(_1531_),
    .S0(net198),
    .S1(net193),
    .X(_3373_));
 sky130_fd_sc_hd__mux2_1 _6429_ (.A0(_3310_),
    .A1(_3373_),
    .S(net205),
    .X(_3374_));
 sky130_fd_sc_hd__nand2_1 _6430_ (.A(net213),
    .B(_3374_),
    .Y(_3375_));
 sky130_fd_sc_hd__o211a_1 _6431_ (.A1(net213),
    .A2(_3231_),
    .B1(_3375_),
    .C1(net190),
    .X(_3376_));
 sky130_fd_sc_hd__a21oi_1 _6432_ (.A1(_2853_),
    .A2(_3058_),
    .B1(_3376_),
    .Y(_3377_));
 sky130_fd_sc_hd__a221o_1 _6433_ (.A1(_1575_),
    .A2(net361),
    .B1(net358),
    .B2(_1578_),
    .C1(net363),
    .X(_3378_));
 sky130_fd_sc_hd__a221o_1 _6434_ (.A1(net189),
    .A2(_3069_),
    .B1(_3378_),
    .B2(_1579_),
    .C1(net223),
    .X(_3379_));
 sky130_fd_sc_hd__a21o_1 _6435_ (.A1(net189),
    .A2(_3063_),
    .B1(_3257_),
    .X(_3380_));
 sky130_fd_sc_hd__o21ai_1 _6436_ (.A1(net319),
    .A2(_3372_),
    .B1(_3380_),
    .Y(_3381_));
 sky130_fd_sc_hd__a21oi_1 _6437_ (.A1(_1578_),
    .A2(net223),
    .B1(net474),
    .Y(_3382_));
 sky130_fd_sc_hd__o31a_2 _6438_ (.A1(_3377_),
    .A2(_3379_),
    .A3(_3381_),
    .B1(_3382_),
    .X(_0836_));
 sky130_fd_sc_hd__xnor2_1 _6439_ (.A(_1599_),
    .B(net359),
    .Y(_3383_));
 sky130_fd_sc_hd__nand2_1 _6440_ (.A(_1601_),
    .B(_3383_),
    .Y(_3384_));
 sky130_fd_sc_hd__nor2_1 _6441_ (.A(_1601_),
    .B(_3383_),
    .Y(_3385_));
 sky130_fd_sc_hd__or2_1 _6442_ (.A(_1601_),
    .B(_3383_),
    .X(_3386_));
 sky130_fd_sc_hd__nand2_1 _6443_ (.A(_3384_),
    .B(_3386_),
    .Y(_3387_));
 sky130_fd_sc_hd__a21o_1 _6444_ (.A1(_3366_),
    .A2(_3368_),
    .B1(_3369_),
    .X(_3388_));
 sky130_fd_sc_hd__xor2_1 _6445_ (.A(_3387_),
    .B(_3388_),
    .X(_3389_));
 sky130_fd_sc_hd__o21a_1 _6446_ (.A1(net185),
    .A2(_3091_),
    .B1(_3256_),
    .X(_3390_));
 sky130_fd_sc_hd__a221o_1 _6447_ (.A1(_1602_),
    .A2(net363),
    .B1(net361),
    .B2(_1599_),
    .C1(net223),
    .X(_3391_));
 sky130_fd_sc_hd__nor2_1 _6448_ (.A(_2864_),
    .B(_3387_),
    .Y(_3392_));
 sky130_fd_sc_hd__a211o_1 _6449_ (.A1(net189),
    .A2(_3094_),
    .B1(_3391_),
    .C1(_3392_),
    .X(_3393_));
 sky130_fd_sc_hd__mux4_1 _6450_ (.A0(_1567_),
    .A1(_1590_),
    .A2(_1601_),
    .A3(_1577_),
    .S0(net192),
    .S1(net200),
    .X(_3394_));
 sky130_fd_sc_hd__mux2_1 _6451_ (.A0(_3323_),
    .A1(_3394_),
    .S(net205),
    .X(_3395_));
 sky130_fd_sc_hd__mux2_1 _6452_ (.A0(_3252_),
    .A1(_3395_),
    .S(net213),
    .X(_3396_));
 sky130_fd_sc_hd__or2_1 _6453_ (.A(net186),
    .B(_3396_),
    .X(_3397_));
 sky130_fd_sc_hd__nand2_1 _6454_ (.A(net186),
    .B(_3081_),
    .Y(_3398_));
 sky130_fd_sc_hd__a32o_1 _6455_ (.A1(_2850_),
    .A2(_3397_),
    .A3(_3398_),
    .B1(_2862_),
    .B2(_3389_),
    .X(_3399_));
 sky130_fd_sc_hd__a21o_1 _6456_ (.A1(_1599_),
    .A2(net2310),
    .B1(net221),
    .X(_3400_));
 sky130_fd_sc_hd__o311a_1 _6457_ (.A1(_3390_),
    .A2(_3393_),
    .A3(_3399_),
    .B1(net2311),
    .C1(net454),
    .X(_0837_));
 sky130_fd_sc_hd__a21o_1 _6458_ (.A1(_3384_),
    .A2(_3388_),
    .B1(_3385_),
    .X(_3401_));
 sky130_fd_sc_hd__xnor2_1 _6459_ (.A(_1634_),
    .B(net359),
    .Y(_3402_));
 sky130_fd_sc_hd__nand2_1 _6460_ (.A(_1637_),
    .B(_3402_),
    .Y(_3403_));
 sky130_fd_sc_hd__nor2_1 _6461_ (.A(_1637_),
    .B(_3402_),
    .Y(_3404_));
 sky130_fd_sc_hd__inv_2 _6462_ (.A(_3404_),
    .Y(_3405_));
 sky130_fd_sc_hd__nand2_1 _6463_ (.A(_3403_),
    .B(_3405_),
    .Y(_3406_));
 sky130_fd_sc_hd__xnor2_1 _6464_ (.A(_3401_),
    .B(_3406_),
    .Y(_3407_));
 sky130_fd_sc_hd__mux4_1 _6465_ (.A0(_1577_),
    .A1(_1637_),
    .A2(_1567_),
    .A3(_1601_),
    .S0(net200),
    .S1(net192),
    .X(_3408_));
 sky130_fd_sc_hd__mux2_1 _6466_ (.A0(_3340_),
    .A1(_3408_),
    .S(net206),
    .X(_3409_));
 sky130_fd_sc_hd__mux2_1 _6467_ (.A0(_3273_),
    .A1(_3409_),
    .S(net214),
    .X(_3410_));
 sky130_fd_sc_hd__nor2_1 _6468_ (.A(net186),
    .B(_3410_),
    .Y(_3411_));
 sky130_fd_sc_hd__a211o_1 _6469_ (.A1(net186),
    .A2(_3107_),
    .B1(_3411_),
    .C1(_2851_),
    .X(_3412_));
 sky130_fd_sc_hd__a21oi_1 _6470_ (.A1(_1634_),
    .A2(net361),
    .B1(net363),
    .Y(_3413_));
 sky130_fd_sc_hd__o21a_1 _6471_ (.A1(_1638_),
    .A2(_2864_),
    .B1(_3413_),
    .X(_3414_));
 sky130_fd_sc_hd__a31o_1 _6472_ (.A1(net189),
    .A2(_3110_),
    .A3(_3111_),
    .B1(_3257_),
    .X(_3415_));
 sky130_fd_sc_hd__o32a_1 _6473_ (.A1(net185),
    .A2(_2819_),
    .A3(_3111_),
    .B1(_3414_),
    .B2(_1639_),
    .X(_3416_));
 sky130_fd_sc_hd__and4_1 _6474_ (.A(net221),
    .B(_3412_),
    .C(_3415_),
    .D(_3416_),
    .X(_3417_));
 sky130_fd_sc_hd__o21a_1 _6475_ (.A1(net319),
    .A2(_3407_),
    .B1(_3417_),
    .X(_3418_));
 sky130_fd_sc_hd__nor2_1 _6476_ (.A(_1638_),
    .B(net221),
    .Y(_3419_));
 sky130_fd_sc_hd__nor3_1 _6477_ (.A(net474),
    .B(_3418_),
    .C(_3419_),
    .Y(_0838_));
 sky130_fd_sc_hd__xnor2_1 _6478_ (.A(_1611_),
    .B(net359),
    .Y(_3420_));
 sky130_fd_sc_hd__and2_1 _6479_ (.A(_1614_),
    .B(_3420_),
    .X(_3421_));
 sky130_fd_sc_hd__nand2_1 _6480_ (.A(_1614_),
    .B(_3420_),
    .Y(_3422_));
 sky130_fd_sc_hd__nor2_1 _6481_ (.A(_1614_),
    .B(_3420_),
    .Y(_3423_));
 sky130_fd_sc_hd__nor2_1 _6482_ (.A(_3421_),
    .B(_3423_),
    .Y(_3424_));
 sky130_fd_sc_hd__a21o_1 _6483_ (.A1(_3401_),
    .A2(_3403_),
    .B1(_3404_),
    .X(_3425_));
 sky130_fd_sc_hd__nand2_1 _6484_ (.A(_3424_),
    .B(_3425_),
    .Y(_3426_));
 sky130_fd_sc_hd__or2_1 _6485_ (.A(_3424_),
    .B(_3425_),
    .X(_3427_));
 sky130_fd_sc_hd__a21oi_1 _6486_ (.A1(_3426_),
    .A2(_3427_),
    .B1(net319),
    .Y(_3428_));
 sky130_fd_sc_hd__mux4_1 _6487_ (.A0(_1601_),
    .A1(_1614_),
    .A2(_1577_),
    .A3(_1637_),
    .S0(net200),
    .S1(net192),
    .X(_3429_));
 sky130_fd_sc_hd__mux2_1 _6488_ (.A0(_3360_),
    .A1(_3429_),
    .S(net206),
    .X(_3430_));
 sky130_fd_sc_hd__mux2_1 _6489_ (.A0(_3289_),
    .A1(_3430_),
    .S(net213),
    .X(_3431_));
 sky130_fd_sc_hd__o2bb2a_1 _6490_ (.A1_N(_2853_),
    .A2_N(_3129_),
    .B1(_3431_),
    .B2(net186),
    .X(_3432_));
 sky130_fd_sc_hd__a21oi_1 _6491_ (.A1(net189),
    .A2(_3135_),
    .B1(_3257_),
    .Y(_3433_));
 sky130_fd_sc_hd__a221o_1 _6492_ (.A1(_1615_),
    .A2(net363),
    .B1(net361),
    .B2(_1611_),
    .C1(net223),
    .X(_3434_));
 sky130_fd_sc_hd__a31o_1 _6493_ (.A1(net189),
    .A2(_2884_),
    .A3(_3065_),
    .B1(_3433_),
    .X(_3435_));
 sky130_fd_sc_hd__a211o_1 _6494_ (.A1(net358),
    .A2(_3424_),
    .B1(_3434_),
    .C1(_3435_),
    .X(_3436_));
 sky130_fd_sc_hd__a21o_1 _6495_ (.A1(_1611_),
    .A2(_1614_),
    .B1(net221),
    .X(_3437_));
 sky130_fd_sc_hd__o311a_1 _6496_ (.A1(_3428_),
    .A2(_3432_),
    .A3(_3436_),
    .B1(_3437_),
    .C1(net446),
    .X(_0839_));
 sky130_fd_sc_hd__a21o_1 _6497_ (.A1(_3422_),
    .A2(_3425_),
    .B1(_3423_),
    .X(_3438_));
 sky130_fd_sc_hd__xnor2_1 _6498_ (.A(_1622_),
    .B(net359),
    .Y(_3439_));
 sky130_fd_sc_hd__nor2_1 _6499_ (.A(_1624_),
    .B(_3439_),
    .Y(_3440_));
 sky130_fd_sc_hd__nand2_1 _6500_ (.A(_1624_),
    .B(_3439_),
    .Y(_3441_));
 sky130_fd_sc_hd__and2b_1 _6501_ (.A_N(_3440_),
    .B(_3441_),
    .X(_3442_));
 sky130_fd_sc_hd__xnor2_1 _6502_ (.A(_3438_),
    .B(_3442_),
    .Y(_3443_));
 sky130_fd_sc_hd__mux4_1 _6503_ (.A0(_1624_),
    .A1(_1637_),
    .A2(_1614_),
    .A3(_1601_),
    .S0(net197),
    .S1(net194),
    .X(_3444_));
 sky130_fd_sc_hd__mux2_1 _6504_ (.A0(_3373_),
    .A1(_3444_),
    .S(net205),
    .X(_3445_));
 sky130_fd_sc_hd__mux2_1 _6505_ (.A0(_3311_),
    .A1(_3445_),
    .S(net213),
    .X(_3446_));
 sky130_fd_sc_hd__o2bb2a_1 _6506_ (.A1_N(_2853_),
    .A2_N(_3150_),
    .B1(_3446_),
    .B2(net186),
    .X(_3447_));
 sky130_fd_sc_hd__a21oi_1 _6507_ (.A1(net189),
    .A2(_3156_),
    .B1(_3257_),
    .Y(_3448_));
 sky130_fd_sc_hd__a2bb2o_1 _6508_ (.A1_N(_2864_),
    .A2_N(_1625_),
    .B1(_1622_),
    .B2(net361),
    .X(_3449_));
 sky130_fd_sc_hd__o21ba_1 _6509_ (.A1(net363),
    .A2(_3449_),
    .B1_N(_1626_),
    .X(_3450_));
 sky130_fd_sc_hd__a311o_1 _6510_ (.A1(net189),
    .A2(_2929_),
    .A3(_3065_),
    .B1(_3450_),
    .C1(net223),
    .X(_3451_));
 sky130_fd_sc_hd__a211o_1 _6511_ (.A1(_2862_),
    .A2(_3443_),
    .B1(_3447_),
    .C1(_3451_),
    .X(_3452_));
 sky130_fd_sc_hd__o221a_1 _6512_ (.A1(_1625_),
    .A2(net221),
    .B1(_3448_),
    .B2(_3452_),
    .C1(net454),
    .X(_0840_));
 sky130_fd_sc_hd__xnor2_1 _6513_ (.A(_1647_),
    .B(net359),
    .Y(_3453_));
 sky130_fd_sc_hd__nor2_1 _6514_ (.A(_1649_),
    .B(_3453_),
    .Y(_3454_));
 sky130_fd_sc_hd__nand2_1 _6515_ (.A(_1649_),
    .B(_3453_),
    .Y(_3455_));
 sky130_fd_sc_hd__nand2b_1 _6516_ (.A_N(_3454_),
    .B(_3455_),
    .Y(_3456_));
 sky130_fd_sc_hd__a21o_1 _6517_ (.A1(_3438_),
    .A2(_3441_),
    .B1(_3440_),
    .X(_3457_));
 sky130_fd_sc_hd__xor2_1 _6518_ (.A(_3456_),
    .B(_3457_),
    .X(_3458_));
 sky130_fd_sc_hd__nand2_1 _6519_ (.A(_2862_),
    .B(_3458_),
    .Y(_3459_));
 sky130_fd_sc_hd__mux4_1 _6520_ (.A0(_1614_),
    .A1(_1637_),
    .A2(_1649_),
    .A3(_1624_),
    .S0(net194),
    .S1(net200),
    .X(_3460_));
 sky130_fd_sc_hd__mux2_1 _6521_ (.A0(_3394_),
    .A1(_3460_),
    .S(net205),
    .X(_3461_));
 sky130_fd_sc_hd__mux2_1 _6522_ (.A0(_3324_),
    .A1(_3461_),
    .S(net213),
    .X(_3462_));
 sky130_fd_sc_hd__a2bb2o_1 _6523_ (.A1_N(net186),
    .A2_N(_3462_),
    .B1(_3172_),
    .B2(_2853_),
    .X(_3463_));
 sky130_fd_sc_hd__o21ai_1 _6524_ (.A1(net185),
    .A2(_3177_),
    .B1(_3256_),
    .Y(_3464_));
 sky130_fd_sc_hd__a21o_1 _6525_ (.A1(_1647_),
    .A2(net361),
    .B1(net363),
    .X(_3465_));
 sky130_fd_sc_hd__o21ai_1 _6526_ (.A1(_1647_),
    .A2(_1649_),
    .B1(_3465_),
    .Y(_3466_));
 sky130_fd_sc_hd__o211a_1 _6527_ (.A1(_2864_),
    .A2(_3456_),
    .B1(_3466_),
    .C1(net221),
    .X(_3467_));
 sky130_fd_sc_hd__o311a_1 _6528_ (.A1(net185),
    .A2(_2959_),
    .A3(_3066_),
    .B1(_3464_),
    .C1(_3467_),
    .X(_3468_));
 sky130_fd_sc_hd__a21oi_1 _6529_ (.A1(_1647_),
    .A2(_1649_),
    .B1(net221),
    .Y(_3469_));
 sky130_fd_sc_hd__a311oi_1 _6530_ (.A1(_3459_),
    .A2(_3463_),
    .A3(_3468_),
    .B1(_3469_),
    .C1(net474),
    .Y(_0841_));
 sky130_fd_sc_hd__a21o_1 _6531_ (.A1(_3455_),
    .A2(_3457_),
    .B1(_3454_),
    .X(_3470_));
 sky130_fd_sc_hd__xnor2_1 _6532_ (.A(_1477_),
    .B(net359),
    .Y(_3471_));
 sky130_fd_sc_hd__nor2_1 _6533_ (.A(_1480_),
    .B(_3471_),
    .Y(_3472_));
 sky130_fd_sc_hd__nand2_1 _6534_ (.A(_1480_),
    .B(_3471_),
    .Y(_3473_));
 sky130_fd_sc_hd__nand2b_1 _6535_ (.A_N(_3472_),
    .B(_3473_),
    .Y(_3474_));
 sky130_fd_sc_hd__xnor2_1 _6536_ (.A(_3470_),
    .B(_3474_),
    .Y(_3475_));
 sky130_fd_sc_hd__nor2_1 _6537_ (.A(net319),
    .B(_3475_),
    .Y(_3476_));
 sky130_fd_sc_hd__mux4_1 _6538_ (.A0(_1480_),
    .A1(_1624_),
    .A2(_1649_),
    .A3(_1614_),
    .S0(net197),
    .S1(net192),
    .X(_3477_));
 sky130_fd_sc_hd__mux2_1 _6539_ (.A0(_3408_),
    .A1(_3477_),
    .S(net206),
    .X(_3478_));
 sky130_fd_sc_hd__mux2_1 _6540_ (.A0(_3341_),
    .A1(_3478_),
    .S(net214),
    .X(_3479_));
 sky130_fd_sc_hd__o22a_1 _6541_ (.A1(_2852_),
    .A2(_3192_),
    .B1(_3479_),
    .B2(net187),
    .X(_3480_));
 sky130_fd_sc_hd__o21a_1 _6542_ (.A1(net185),
    .A2(_3198_),
    .B1(_3256_),
    .X(_3481_));
 sky130_fd_sc_hd__a221o_1 _6543_ (.A1(_1477_),
    .A2(net361),
    .B1(net358),
    .B2(_1481_),
    .C1(net363),
    .X(_3482_));
 sky130_fd_sc_hd__a21o_1 _6544_ (.A1(_1482_),
    .A2(_3482_),
    .B1(net223),
    .X(_3483_));
 sky130_fd_sc_hd__a311o_1 _6545_ (.A1(net212),
    .A2(_2996_),
    .A3(_3276_),
    .B1(_3481_),
    .C1(_3483_),
    .X(_3484_));
 sky130_fd_sc_hd__nand2_1 _6546_ (.A(_1481_),
    .B(net223),
    .Y(_3485_));
 sky130_fd_sc_hd__o311a_1 _6547_ (.A1(_3476_),
    .A2(_3480_),
    .A3(_3484_),
    .B1(_3485_),
    .C1(net446),
    .X(_0842_));
 sky130_fd_sc_hd__xnor2_1 _6548_ (.A(_1500_),
    .B(net359),
    .Y(_3486_));
 sky130_fd_sc_hd__nor2_1 _6549_ (.A(_1503_),
    .B(_3486_),
    .Y(_3487_));
 sky130_fd_sc_hd__nand2_1 _6550_ (.A(_1503_),
    .B(_3486_),
    .Y(_3488_));
 sky130_fd_sc_hd__nand2b_1 _6551_ (.A_N(_3487_),
    .B(_3488_),
    .Y(_3489_));
 sky130_fd_sc_hd__a21o_1 _6552_ (.A1(_3470_),
    .A2(_3473_),
    .B1(_3472_),
    .X(_3490_));
 sky130_fd_sc_hd__xnor2_1 _6553_ (.A(_3489_),
    .B(_3490_),
    .Y(_3491_));
 sky130_fd_sc_hd__mux4_1 _6554_ (.A0(_1503_),
    .A1(_1649_),
    .A2(_1480_),
    .A3(_1624_),
    .S0(net197),
    .S1(net194),
    .X(_3492_));
 sky130_fd_sc_hd__mux2_1 _6555_ (.A0(_3429_),
    .A1(_3492_),
    .S(net205),
    .X(_3493_));
 sky130_fd_sc_hd__mux2_1 _6556_ (.A0(_3361_),
    .A1(_3493_),
    .S(net214),
    .X(_3494_));
 sky130_fd_sc_hd__a2bb2o_1 _6557_ (.A1_N(net187),
    .A2_N(_3494_),
    .B1(_3211_),
    .B2(_2853_),
    .X(_3495_));
 sky130_fd_sc_hd__a21o_1 _6558_ (.A1(net189),
    .A2(_3217_),
    .B1(_3257_),
    .X(_3496_));
 sky130_fd_sc_hd__a221o_1 _6559_ (.A1(_1504_),
    .A2(net363),
    .B1(net361),
    .B2(_1500_),
    .C1(net223),
    .X(_3497_));
 sky130_fd_sc_hd__o21ba_1 _6560_ (.A1(_2864_),
    .A2(_3489_),
    .B1_N(_3497_),
    .X(_3498_));
 sky130_fd_sc_hd__o311a_1 _6561_ (.A1(net185),
    .A2(_3025_),
    .A3(_3066_),
    .B1(_3496_),
    .C1(_3498_),
    .X(_3499_));
 sky130_fd_sc_hd__o211a_1 _6562_ (.A1(net319),
    .A2(_3491_),
    .B1(_3495_),
    .C1(_3499_),
    .X(_3500_));
 sky130_fd_sc_hd__a21oi_1 _6563_ (.A1(net2299),
    .A2(_1503_),
    .B1(net221),
    .Y(_3501_));
 sky130_fd_sc_hd__nor3_1 _6564_ (.A(net475),
    .B(_3500_),
    .C(net2300),
    .Y(_0843_));
 sky130_fd_sc_hd__a21o_1 _6565_ (.A1(_3488_),
    .A2(_3490_),
    .B1(_3487_),
    .X(_3502_));
 sky130_fd_sc_hd__xnor2_1 _6566_ (.A(_1488_),
    .B(_2859_),
    .Y(_3503_));
 sky130_fd_sc_hd__inv_2 _6567_ (.A(_3503_),
    .Y(_3504_));
 sky130_fd_sc_hd__nor2_1 _6568_ (.A(_1490_),
    .B(_3504_),
    .Y(_3505_));
 sky130_fd_sc_hd__nand2_1 _6569_ (.A(_1490_),
    .B(_3504_),
    .Y(_3506_));
 sky130_fd_sc_hd__nand2b_1 _6570_ (.A_N(_3505_),
    .B(_3506_),
    .Y(_3507_));
 sky130_fd_sc_hd__xnor2_1 _6571_ (.A(_3502_),
    .B(_3507_),
    .Y(_3508_));
 sky130_fd_sc_hd__mux4_1 _6572_ (.A0(_1480_),
    .A1(_1490_),
    .A2(_1649_),
    .A3(_1503_),
    .S0(net200),
    .S1(net192),
    .X(_3509_));
 sky130_fd_sc_hd__mux2_1 _6573_ (.A0(_3444_),
    .A1(_3509_),
    .S(net205),
    .X(_3510_));
 sky130_fd_sc_hd__mux2_1 _6574_ (.A0(_3374_),
    .A1(_3510_),
    .S(net213),
    .X(_3511_));
 sky130_fd_sc_hd__a2bb2o_1 _6575_ (.A1_N(net186),
    .A2_N(_3511_),
    .B1(_3233_),
    .B2(_2853_),
    .X(_3512_));
 sky130_fd_sc_hd__o21ai_1 _6576_ (.A1(net185),
    .A2(_3238_),
    .B1(_3256_),
    .Y(_3513_));
 sky130_fd_sc_hd__a221o_1 _6577_ (.A1(_1488_),
    .A2(net361),
    .B1(net358),
    .B2(_1491_),
    .C1(net363),
    .X(_3514_));
 sky130_fd_sc_hd__o21ai_1 _6578_ (.A1(_1488_),
    .A2(_1490_),
    .B1(_3514_),
    .Y(_3515_));
 sky130_fd_sc_hd__o311a_1 _6579_ (.A1(net185),
    .A2(_3066_),
    .A3(_3067_),
    .B1(_3515_),
    .C1(net221),
    .X(_3516_));
 sky130_fd_sc_hd__o211a_1 _6580_ (.A1(net319),
    .A2(_3508_),
    .B1(_3513_),
    .C1(_3516_),
    .X(_3517_));
 sky130_fd_sc_hd__a221oi_1 _6581_ (.A1(_1491_),
    .A2(net223),
    .B1(_3512_),
    .B2(_3517_),
    .C1(net475),
    .Y(_0844_));
 sky130_fd_sc_hd__a21oi_1 _6582_ (.A1(_3502_),
    .A2(_3506_),
    .B1(_3505_),
    .Y(_3518_));
 sky130_fd_sc_hd__and2_1 _6583_ (.A(_1469_),
    .B(net359),
    .X(_3519_));
 sky130_fd_sc_hd__nor2_1 _6584_ (.A(_1469_),
    .B(net359),
    .Y(_3520_));
 sky130_fd_sc_hd__nor2_1 _6585_ (.A(_3519_),
    .B(_3520_),
    .Y(_3521_));
 sky130_fd_sc_hd__a211o_1 _6586_ (.A1(_3502_),
    .A2(_3506_),
    .B1(_3521_),
    .C1(_3505_),
    .X(_3522_));
 sky130_fd_sc_hd__o311a_1 _6587_ (.A1(_3518_),
    .A2(_3519_),
    .A3(_3520_),
    .B1(_3522_),
    .C1(_2862_),
    .X(_3523_));
 sky130_fd_sc_hd__mux4_1 _6588_ (.A0(_1467_),
    .A1(_1490_),
    .A2(_1503_),
    .A3(_1480_),
    .S0(net192),
    .S1(net197),
    .X(_3524_));
 sky130_fd_sc_hd__or2_1 _6589_ (.A(net202),
    .B(_3524_),
    .X(_3525_));
 sky130_fd_sc_hd__o211a_1 _6590_ (.A1(net205),
    .A2(_3460_),
    .B1(_3525_),
    .C1(net212),
    .X(_3526_));
 sky130_fd_sc_hd__a211o_1 _6591_ (.A1(net208),
    .A2(_3395_),
    .B1(_3526_),
    .C1(net186),
    .X(_3527_));
 sky130_fd_sc_hd__o211a_1 _6592_ (.A1(net190),
    .A2(_3253_),
    .B1(_3527_),
    .C1(_2850_),
    .X(_3528_));
 sky130_fd_sc_hd__o21a_1 _6593_ (.A1(_1451_),
    .A2(_1467_),
    .B1(net363),
    .X(_3529_));
 sky130_fd_sc_hd__a221o_1 _6594_ (.A1(_1467_),
    .A2(_2816_),
    .B1(net361),
    .B2(_1451_),
    .C1(net223),
    .X(_3530_));
 sky130_fd_sc_hd__a211o_1 _6595_ (.A1(_1469_),
    .A2(net358),
    .B1(_3529_),
    .C1(_3530_),
    .X(_3531_));
 sky130_fd_sc_hd__a31o_1 _6596_ (.A1(net212),
    .A2(_3093_),
    .A3(_3276_),
    .B1(_3531_),
    .X(_3532_));
 sky130_fd_sc_hd__a21o_1 _6597_ (.A1(_1451_),
    .A2(_1467_),
    .B1(net221),
    .X(_3533_));
 sky130_fd_sc_hd__o311a_1 _6598_ (.A1(_3523_),
    .A2(_3528_),
    .A3(_3532_),
    .B1(_3533_),
    .C1(net454),
    .X(_0845_));
 sky130_fd_sc_hd__and2_1 _6599_ (.A(net449),
    .B(net2031),
    .X(_0846_));
 sky130_fd_sc_hd__and2_1 _6600_ (.A(net459),
    .B(net1435),
    .X(_0847_));
 sky130_fd_sc_hd__and2_1 _6601_ (.A(net464),
    .B(net1939),
    .X(_0848_));
 sky130_fd_sc_hd__and2_2 _6602_ (.A(net452),
    .B(_1697_),
    .X(_0849_));
 sky130_fd_sc_hd__o31a_4 _6603_ (.A1(_1680_),
    .A2(_1681_),
    .A3(_1682_),
    .B1(net461),
    .X(_0850_));
 sky130_fd_sc_hd__and2_1 _6604_ (.A(net448),
    .B(_1669_),
    .X(_0851_));
 sky130_fd_sc_hd__nor2_1 _6605_ (.A(net480),
    .B(net2121),
    .Y(_0852_));
 sky130_fd_sc_hd__and2_1 _6606_ (.A(net469),
    .B(_1718_),
    .X(_0853_));
 sky130_fd_sc_hd__o31a_1 _6607_ (.A1(_1742_),
    .A2(_1743_),
    .A3(_1744_),
    .B1(net458),
    .X(_0854_));
 sky130_fd_sc_hd__and2_1 _6608_ (.A(net455),
    .B(net2176),
    .X(_0855_));
 sky130_fd_sc_hd__and2_1 _6609_ (.A(net444),
    .B(_1709_),
    .X(_0856_));
 sky130_fd_sc_hd__nor2_1 _6610_ (.A(net475),
    .B(_1779_),
    .Y(_0857_));
 sky130_fd_sc_hd__and2_1 _6611_ (.A(net457),
    .B(_1759_),
    .X(_0858_));
 sky130_fd_sc_hd__and2_1 _6612_ (.A(net469),
    .B(net2174),
    .X(_0859_));
 sky130_fd_sc_hd__and2_1 _6613_ (.A(net440),
    .B(_1790_),
    .X(_0860_));
 sky130_fd_sc_hd__nor2_1 _6614_ (.A(net478),
    .B(_1823_),
    .Y(_0861_));
 sky130_fd_sc_hd__and2_1 _6615_ (.A(net444),
    .B(_1802_),
    .X(_0862_));
 sky130_fd_sc_hd__and2_1 _6616_ (.A(net455),
    .B(_1812_),
    .X(_0863_));
 sky130_fd_sc_hd__and2_1 _6617_ (.A(net457),
    .B(_1836_),
    .X(_0864_));
 sky130_fd_sc_hd__nor2_1 _6618_ (.A(net478),
    .B(net618),
    .Y(_0865_));
 sky130_fd_sc_hd__a31oi_2 _6619_ (.A1(_1513_),
    .A2(_1514_),
    .A3(_1515_),
    .B1(net477),
    .Y(_0866_));
 sky130_fd_sc_hd__and2_1 _6620_ (.A(net465),
    .B(_1552_),
    .X(_0867_));
 sky130_fd_sc_hd__and2_1 _6621_ (.A(net455),
    .B(_1528_),
    .X(_0868_));
 sky130_fd_sc_hd__nor2_1 _6622_ (.A(net475),
    .B(net2141),
    .Y(_0869_));
 sky130_fd_sc_hd__and2_1 _6623_ (.A(net441),
    .B(net2304),
    .X(_0870_));
 sky130_fd_sc_hd__and2_1 _6624_ (.A(net466),
    .B(_1574_),
    .X(_0871_));
 sky130_fd_sc_hd__nor2_1 _6625_ (.A(net473),
    .B(_1597_),
    .Y(_0872_));
 sky130_fd_sc_hd__nor2_1 _6626_ (.A(net481),
    .B(_1632_),
    .Y(_0873_));
 sky130_fd_sc_hd__nor2_1 _6627_ (.A(net474),
    .B(_1609_),
    .Y(_0874_));
 sky130_fd_sc_hd__and2_1 _6628_ (.A(net441),
    .B(_1621_),
    .X(_0875_));
 sky130_fd_sc_hd__nor2_2 _6629_ (.A(net477),
    .B(_1645_),
    .Y(_0876_));
 sky130_fd_sc_hd__nor2_1 _6630_ (.A(net475),
    .B(_1475_),
    .Y(_0877_));
 sky130_fd_sc_hd__nor2_1 _6631_ (.A(net475),
    .B(_1498_),
    .Y(_0878_));
 sky130_fd_sc_hd__and2_1 _6632_ (.A(net450),
    .B(_1487_),
    .X(_0879_));
 sky130_fd_sc_hd__nor2_2 _6633_ (.A(net474),
    .B(_1449_),
    .Y(_0880_));
 sky130_fd_sc_hd__and2_1 _6634_ (.A(net449),
    .B(net841),
    .X(_0881_));
 sky130_fd_sc_hd__and2_1 _6635_ (.A(net465),
    .B(net739),
    .X(_0882_));
 sky130_fd_sc_hd__and2_1 _6636_ (.A(net469),
    .B(net621),
    .X(_0883_));
 sky130_fd_sc_hd__and2_1 _6637_ (.A(net447),
    .B(net849),
    .X(_0884_));
 sky130_fd_sc_hd__and2_1 _6638_ (.A(net469),
    .B(net731),
    .X(_0885_));
 sky130_fd_sc_hd__mux2_1 _6639_ (.A0(net2118),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .S(net481),
    .X(_0886_));
 sky130_fd_sc_hd__mux2_1 _6640_ (.A0(net2039),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .S(net481),
    .X(_0887_));
 sky130_fd_sc_hd__mux2_1 _6641_ (.A0(net2100),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .S(net481),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _6642_ (.A0(net2112),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .S(net481),
    .X(_0889_));
 sky130_fd_sc_hd__and2_1 _6643_ (.A(net470),
    .B(net741),
    .X(_0890_));
 sky130_fd_sc_hd__and2_1 _6644_ (.A(net464),
    .B(net751),
    .X(_0891_));
 sky130_fd_sc_hd__and2_1 _6645_ (.A(net466),
    .B(net723),
    .X(_0892_));
 sky130_fd_sc_hd__and2_1 _6646_ (.A(net456),
    .B(net737),
    .X(_0893_));
 sky130_fd_sc_hd__and2_1 _6647_ (.A(net460),
    .B(net825),
    .X(_0894_));
 sky130_fd_sc_hd__and2_1 _6648_ (.A(net456),
    .B(net745),
    .X(_0895_));
 sky130_fd_sc_hd__and2_1 _6649_ (.A(net455),
    .B(net717),
    .X(_0896_));
 sky130_fd_sc_hd__and2_1 _6650_ (.A(net459),
    .B(net687),
    .X(_0897_));
 sky130_fd_sc_hd__and2_1 _6651_ (.A(net449),
    .B(net659),
    .X(_0898_));
 sky130_fd_sc_hd__and2_1 _6652_ (.A(net447),
    .B(net757),
    .X(_0899_));
 sky130_fd_sc_hd__and2_1 _6653_ (.A(net449),
    .B(net619),
    .X(_0900_));
 sky130_fd_sc_hd__and2_1 _6654_ (.A(net456),
    .B(net781),
    .X(_0901_));
 sky130_fd_sc_hd__and2_1 _6655_ (.A(net457),
    .B(net629),
    .X(_0902_));
 sky130_fd_sc_hd__and2_1 _6656_ (.A(net457),
    .B(net779),
    .X(_0903_));
 sky130_fd_sc_hd__and2_1 _6657_ (.A(net462),
    .B(net695),
    .X(_0904_));
 sky130_fd_sc_hd__and2_1 _6658_ (.A(net457),
    .B(net785),
    .X(_0905_));
 sky130_fd_sc_hd__and2_1 _6659_ (.A(net465),
    .B(net711),
    .X(_0906_));
 sky130_fd_sc_hd__and2_1 _6660_ (.A(net458),
    .B(net809),
    .X(_0907_));
 sky130_fd_sc_hd__and2_1 _6661_ (.A(net470),
    .B(net765),
    .X(_0908_));
 sky130_fd_sc_hd__and2_1 _6662_ (.A(net450),
    .B(net691),
    .X(_0909_));
 sky130_fd_sc_hd__and2_1 _6663_ (.A(net451),
    .B(net635),
    .X(_0910_));
 sky130_fd_sc_hd__and2_1 _6664_ (.A(net450),
    .B(net683),
    .X(_0911_));
 sky130_fd_sc_hd__and2_1 _6665_ (.A(net452),
    .B(net653),
    .X(_0912_));
 sky130_fd_sc_hd__and2_1 _6666_ (.A(net445),
    .B(net829),
    .X(_0913_));
 sky130_fd_sc_hd__and2_1 _6667_ (.A(net445),
    .B(net777),
    .X(_0914_));
 sky130_fd_sc_hd__and2_1 _6668_ (.A(net451),
    .B(net839),
    .X(_0915_));
 sky130_fd_sc_hd__and2_1 _6669_ (.A(net441),
    .B(net645),
    .X(_0916_));
 sky130_fd_sc_hd__and2_1 _6670_ (.A(net447),
    .B(net805),
    .X(_0917_));
 sky130_fd_sc_hd__and2_1 _6671_ (.A(net447),
    .B(net707),
    .X(_0918_));
 sky130_fd_sc_hd__and2_1 _6672_ (.A(net451),
    .B(net697),
    .X(_0919_));
 sky130_fd_sc_hd__and2_1 _6673_ (.A(net462),
    .B(net795),
    .X(_0920_));
 sky130_fd_sc_hd__and2_1 _6674_ (.A(net460),
    .B(net799),
    .X(_0921_));
 sky130_fd_sc_hd__and2_1 _6675_ (.A(net470),
    .B(net771),
    .X(_0922_));
 sky130_fd_sc_hd__and2_1 _6676_ (.A(net464),
    .B(net797),
    .X(_0923_));
 sky130_fd_sc_hd__and2_1 _6677_ (.A(net466),
    .B(net729),
    .X(_0924_));
 sky130_fd_sc_hd__and2_1 _6678_ (.A(net456),
    .B(net759),
    .X(_0925_));
 sky130_fd_sc_hd__and2_1 _6679_ (.A(net460),
    .B(net783),
    .X(_0926_));
 sky130_fd_sc_hd__and2_1 _6680_ (.A(net459),
    .B(net705),
    .X(_0927_));
 sky130_fd_sc_hd__and2_1 _6681_ (.A(net455),
    .B(net709),
    .X(_0928_));
 sky130_fd_sc_hd__and2_1 _6682_ (.A(net459),
    .B(net827),
    .X(_0929_));
 sky130_fd_sc_hd__and2_1 _6683_ (.A(net449),
    .B(net665),
    .X(_0930_));
 sky130_fd_sc_hd__and2_1 _6684_ (.A(net447),
    .B(net669),
    .X(_0931_));
 sky130_fd_sc_hd__and2_1 _6685_ (.A(net455),
    .B(net703),
    .X(_0932_));
 sky130_fd_sc_hd__and2_1 _6686_ (.A(net456),
    .B(net833),
    .X(_0933_));
 sky130_fd_sc_hd__and2_1 _6687_ (.A(net457),
    .B(net819),
    .X(_0934_));
 sky130_fd_sc_hd__and2_1 _6688_ (.A(net457),
    .B(net631),
    .X(_0935_));
 sky130_fd_sc_hd__and2_1 _6689_ (.A(net462),
    .B(net719),
    .X(_0936_));
 sky130_fd_sc_hd__and2_1 _6690_ (.A(net458),
    .B(net831),
    .X(_0937_));
 sky130_fd_sc_hd__and2_1 _6691_ (.A(net465),
    .B(net721),
    .X(_0938_));
 sky130_fd_sc_hd__and2_1 _6692_ (.A(net458),
    .B(net787),
    .X(_0939_));
 sky130_fd_sc_hd__and2_1 _6693_ (.A(net469),
    .B(net647),
    .X(_0940_));
 sky130_fd_sc_hd__and2_1 _6694_ (.A(net450),
    .B(net813),
    .X(_0941_));
 sky130_fd_sc_hd__and2_1 _6695_ (.A(net450),
    .B(net725),
    .X(_0942_));
 sky130_fd_sc_hd__and2_1 _6696_ (.A(net450),
    .B(net677),
    .X(_0943_));
 sky130_fd_sc_hd__and2_1 _6697_ (.A(net453),
    .B(net651),
    .X(_0944_));
 sky130_fd_sc_hd__and2_1 _6698_ (.A(net445),
    .B(net815),
    .X(_0945_));
 sky130_fd_sc_hd__and2_1 _6699_ (.A(net445),
    .B(net639),
    .X(_0946_));
 sky130_fd_sc_hd__and2_1 _6700_ (.A(net450),
    .B(net847),
    .X(_0947_));
 sky130_fd_sc_hd__and2_1 _6701_ (.A(net441),
    .B(net655),
    .X(_0948_));
 sky130_fd_sc_hd__and2_1 _6702_ (.A(net441),
    .B(net837),
    .X(_0949_));
 sky130_fd_sc_hd__and2_1 _6703_ (.A(net448),
    .B(net675),
    .X(_0950_));
 sky130_fd_sc_hd__and2_1 _6704_ (.A(net451),
    .B(net679),
    .X(_0951_));
 sky130_fd_sc_hd__and2_1 _6705_ (.A(net462),
    .B(net31),
    .X(_0952_));
 sky130_fd_sc_hd__and2_1 _6706_ (.A(net452),
    .B(net42),
    .X(_0953_));
 sky130_fd_sc_hd__and2_1 _6707_ (.A(net470),
    .B(net53),
    .X(_0954_));
 sky130_fd_sc_hd__and2_1 _6708_ (.A(net464),
    .B(net56),
    .X(_0955_));
 sky130_fd_sc_hd__and2_1 _6709_ (.A(net466),
    .B(net57),
    .X(_0956_));
 sky130_fd_sc_hd__and2_1 _6710_ (.A(net455),
    .B(net58),
    .X(_0957_));
 sky130_fd_sc_hd__and2_1 _6711_ (.A(net460),
    .B(net59),
    .X(_0958_));
 sky130_fd_sc_hd__and2_1 _6712_ (.A(net465),
    .B(net60),
    .X(_0959_));
 sky130_fd_sc_hd__and2_1 _6713_ (.A(net455),
    .B(net61),
    .X(_0960_));
 sky130_fd_sc_hd__and2_1 _6714_ (.A(net469),
    .B(net62),
    .X(_0961_));
 sky130_fd_sc_hd__and2_1 _6715_ (.A(net448),
    .B(net32),
    .X(_0962_));
 sky130_fd_sc_hd__and2_1 _6716_ (.A(net440),
    .B(net33),
    .X(_0963_));
 sky130_fd_sc_hd__and2_1 _6717_ (.A(net455),
    .B(net34),
    .X(_0964_));
 sky130_fd_sc_hd__and2_1 _6718_ (.A(net460),
    .B(net35),
    .X(_0965_));
 sky130_fd_sc_hd__and2_1 _6719_ (.A(net449),
    .B(net36),
    .X(_0966_));
 sky130_fd_sc_hd__and2_1 _6720_ (.A(net447),
    .B(net37),
    .X(_0967_));
 sky130_fd_sc_hd__and2_1 _6721_ (.A(net461),
    .B(net38),
    .X(_0968_));
 sky130_fd_sc_hd__and2_1 _6722_ (.A(net466),
    .B(net39),
    .X(_0969_));
 sky130_fd_sc_hd__and2_1 _6723_ (.A(net471),
    .B(net40),
    .X(_0970_));
 sky130_fd_sc_hd__and2_1 _6724_ (.A(net440),
    .B(net41),
    .X(_0971_));
 sky130_fd_sc_hd__and2_1 _6725_ (.A(net470),
    .B(net43),
    .X(_0972_));
 sky130_fd_sc_hd__and2_1 _6726_ (.A(net463),
    .B(net44),
    .X(_0973_));
 sky130_fd_sc_hd__and2_1 _6727_ (.A(net448),
    .B(net45),
    .X(_0974_));
 sky130_fd_sc_hd__and2_1 _6728_ (.A(net450),
    .B(net46),
    .X(_0975_));
 sky130_fd_sc_hd__and2_1 _6729_ (.A(net464),
    .B(net47),
    .X(_0976_));
 sky130_fd_sc_hd__and2_1 _6730_ (.A(net444),
    .B(net48),
    .X(_0977_));
 sky130_fd_sc_hd__and2_1 _6731_ (.A(net445),
    .B(net49),
    .X(_0978_));
 sky130_fd_sc_hd__and2_1 _6732_ (.A(net452),
    .B(net50),
    .X(_0979_));
 sky130_fd_sc_hd__and2_1 _6733_ (.A(net441),
    .B(net51),
    .X(_0980_));
 sky130_fd_sc_hd__and2_1 _6734_ (.A(net449),
    .B(net52),
    .X(_0981_));
 sky130_fd_sc_hd__and2_1 _6735_ (.A(net457),
    .B(net54),
    .X(_0982_));
 sky130_fd_sc_hd__and2_1 _6736_ (.A(net472),
    .B(net55),
    .X(_0983_));
 sky130_fd_sc_hd__and3_1 _6737_ (.A(net2010),
    .B(net179),
    .C(net285),
    .X(_1017_));
 sky130_fd_sc_hd__and3_1 _6738_ (.A(net2092),
    .B(net182),
    .C(net289),
    .X(_1018_));
 sky130_fd_sc_hd__and3_1 _6739_ (.A(net2055),
    .B(net175),
    .C(net279),
    .X(_1019_));
 sky130_fd_sc_hd__nor4_2 _6740_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2744_),
    .D(_2767_),
    .Y(_3534_));
 sky130_fd_sc_hd__inv_2 _6741_ (.A(net316),
    .Y(_3535_));
 sky130_fd_sc_hd__nor2_2 _6742_ (.A(net479),
    .B(net316),
    .Y(_3536_));
 sky130_fd_sc_hd__or2_1 _6743_ (.A(net481),
    .B(net316),
    .X(_3537_));
 sky130_fd_sc_hd__o22a_1 _6744_ (.A1(net331),
    .A2(_3535_),
    .B1(_3537_),
    .B2(net924),
    .X(_1020_));
 sky130_fd_sc_hd__o22a_1 _6745_ (.A1(net332),
    .A2(_3535_),
    .B1(_3537_),
    .B2(net857),
    .X(_1021_));
 sky130_fd_sc_hd__a22o_1 _6746_ (.A1(net333),
    .A2(net316),
    .B1(net259),
    .B2(net1557),
    .X(_1022_));
 sky130_fd_sc_hd__a22o_1 _6747_ (.A1(net334),
    .A2(net316),
    .B1(net259),
    .B2(net1106),
    .X(_1023_));
 sky130_fd_sc_hd__a22o_1 _6748_ (.A1(net329),
    .A2(net318),
    .B1(net259),
    .B2(net1525),
    .X(_1024_));
 sky130_fd_sc_hd__a22o_1 _6749_ (.A1(_1741_),
    .A2(net316),
    .B1(net259),
    .B2(net1637),
    .X(_1025_));
 sky130_fd_sc_hd__a22o_1 _6750_ (.A1(net328),
    .A2(net316),
    .B1(net259),
    .B2(net918),
    .X(_1026_));
 sky130_fd_sc_hd__a22o_1 _6751_ (.A1(net330),
    .A2(net317),
    .B1(net258),
    .B2(net1114),
    .X(_1027_));
 sky130_fd_sc_hd__a22o_1 _6752_ (.A1(net325),
    .A2(net317),
    .B1(net258),
    .B2(net1339),
    .X(_1028_));
 sky130_fd_sc_hd__a22o_1 _6753_ (.A1(net327),
    .A2(net316),
    .B1(net259),
    .B2(net1164),
    .X(_1029_));
 sky130_fd_sc_hd__a22o_1 _6754_ (.A1(net326),
    .A2(net317),
    .B1(net258),
    .B2(net1196),
    .X(_1030_));
 sky130_fd_sc_hd__a22o_1 _6755_ (.A1(net324),
    .A2(net317),
    .B1(net258),
    .B2(net1066),
    .X(_1031_));
 sky130_fd_sc_hd__a22o_1 _6756_ (.A1(net321),
    .A2(net316),
    .B1(net259),
    .B2(net1459),
    .X(_1032_));
 sky130_fd_sc_hd__a22o_1 _6757_ (.A1(net323),
    .A2(net316),
    .B1(net259),
    .B2(net1385),
    .X(_1033_));
 sky130_fd_sc_hd__a22o_1 _6758_ (.A1(net322),
    .A2(net316),
    .B1(net259),
    .B2(net1375),
    .X(_1034_));
 sky130_fd_sc_hd__a22o_1 _6759_ (.A1(net320),
    .A2(net316),
    .B1(net259),
    .B2(net1152),
    .X(_1035_));
 sky130_fd_sc_hd__a22o_1 _6760_ (.A1(net344),
    .A2(net317),
    .B1(net258),
    .B2(net1539),
    .X(_1036_));
 sky130_fd_sc_hd__a22o_1 _6761_ (.A1(_1512_),
    .A2(net317),
    .B1(net258),
    .B2(net1327),
    .X(_1037_));
 sky130_fd_sc_hd__a22o_1 _6762_ (.A1(net343),
    .A2(net316),
    .B1(net259),
    .B2(net952),
    .X(_1038_));
 sky130_fd_sc_hd__a22o_1 _6763_ (.A1(net345),
    .A2(net316),
    .B1(net259),
    .B2(net1347),
    .X(_1039_));
 sky130_fd_sc_hd__a22o_1 _6764_ (.A1(net340),
    .A2(net317),
    .B1(net258),
    .B2(net1098),
    .X(_1040_));
 sky130_fd_sc_hd__a22o_1 _6765_ (.A1(net342),
    .A2(net317),
    .B1(net258),
    .B2(net1276),
    .X(_1041_));
 sky130_fd_sc_hd__a22o_1 _6766_ (.A1(net341),
    .A2(net318),
    .B1(net259),
    .B2(net1232),
    .X(_1042_));
 sky130_fd_sc_hd__a22o_1 _6767_ (.A1(net339),
    .A2(net317),
    .B1(net258),
    .B2(net1515),
    .X(_1043_));
 sky130_fd_sc_hd__a22o_1 _6768_ (.A1(net336),
    .A2(net316),
    .B1(net259),
    .B2(net1728),
    .X(_1044_));
 sky130_fd_sc_hd__a22o_1 _6769_ (.A1(net338),
    .A2(net317),
    .B1(net258),
    .B2(net1044),
    .X(_1045_));
 sky130_fd_sc_hd__a22o_1 _6770_ (.A1(net337),
    .A2(net317),
    .B1(net258),
    .B2(net1038),
    .X(_1046_));
 sky130_fd_sc_hd__a22o_1 _6771_ (.A1(net335),
    .A2(net316),
    .B1(net258),
    .B2(net1589),
    .X(_1047_));
 sky130_fd_sc_hd__a22o_1 _6772_ (.A1(net348),
    .A2(net317),
    .B1(net258),
    .B2(net1058),
    .X(_1048_));
 sky130_fd_sc_hd__a22o_1 _6773_ (.A1(net346),
    .A2(net317),
    .B1(net258),
    .B2(net1343),
    .X(_1049_));
 sky130_fd_sc_hd__a22o_1 _6774_ (.A1(net347),
    .A2(net317),
    .B1(net258),
    .B2(net1425),
    .X(_1050_));
 sky130_fd_sc_hd__a22o_1 _6775_ (.A1(net370),
    .A2(net317),
    .B1(net258),
    .B2(net1593),
    .X(_1051_));
 sky130_fd_sc_hd__or2_4 _6776_ (.A(_1413_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .X(_3538_));
 sky130_fd_sc_hd__nor3_2 _6777_ (.A(_2743_),
    .B(net365),
    .C(_3538_),
    .Y(_3539_));
 sky130_fd_sc_hd__or3_4 _6778_ (.A(_2743_),
    .B(net365),
    .C(_3538_),
    .X(_3540_));
 sky130_fd_sc_hd__and2_1 _6779_ (.A(net331),
    .B(net315),
    .X(_3541_));
 sky130_fd_sc_hd__a31o_1 _6780_ (.A1(net468),
    .A2(net1872),
    .A3(net312),
    .B1(_3541_),
    .X(_1052_));
 sky130_fd_sc_hd__and2_1 _6781_ (.A(net332),
    .B(net315),
    .X(_3542_));
 sky130_fd_sc_hd__a31o_1 _6782_ (.A1(net470),
    .A2(net1768),
    .A3(net312),
    .B1(_3542_),
    .X(_1053_));
 sky130_fd_sc_hd__or3_1 _6783_ (.A(net481),
    .B(net2136),
    .C(net315),
    .X(_3543_));
 sky130_fd_sc_hd__o21a_1 _6784_ (.A1(net333),
    .A2(net312),
    .B1(_3543_),
    .X(_1054_));
 sky130_fd_sc_hd__and2_1 _6785_ (.A(net334),
    .B(net314),
    .X(_3544_));
 sky130_fd_sc_hd__a31o_1 _6786_ (.A1(net467),
    .A2(net1772),
    .A3(net312),
    .B1(_3544_),
    .X(_1055_));
 sky130_fd_sc_hd__and2_1 _6787_ (.A(net329),
    .B(net315),
    .X(_3545_));
 sky130_fd_sc_hd__a31o_1 _6788_ (.A1(net467),
    .A2(net1890),
    .A3(_3540_),
    .B1(_3545_),
    .X(_1056_));
 sky130_fd_sc_hd__nor2_1 _6789_ (.A(_1740_),
    .B(_3540_),
    .Y(_3546_));
 sky130_fd_sc_hd__a31o_1 _6790_ (.A1(net464),
    .A2(net1901),
    .A3(_3540_),
    .B1(_3546_),
    .X(_1057_));
 sky130_fd_sc_hd__and2_1 _6791_ (.A(net328),
    .B(net315),
    .X(_3547_));
 sky130_fd_sc_hd__a31o_1 _6792_ (.A1(net460),
    .A2(net1675),
    .A3(net312),
    .B1(_3547_),
    .X(_1058_));
 sky130_fd_sc_hd__and2_1 _6793_ (.A(net330),
    .B(net314),
    .X(_3548_));
 sky130_fd_sc_hd__a31o_1 _6794_ (.A1(net446),
    .A2(net1972),
    .A3(net313),
    .B1(_3548_),
    .X(_1059_));
 sky130_fd_sc_hd__and2_1 _6795_ (.A(net325),
    .B(net314),
    .X(_3549_));
 sky130_fd_sc_hd__a31o_1 _6796_ (.A1(net448),
    .A2(net1974),
    .A3(net313),
    .B1(_3549_),
    .X(_1060_));
 sky130_fd_sc_hd__and2_1 _6797_ (.A(net327),
    .B(net315),
    .X(_3550_));
 sky130_fd_sc_hd__a31o_1 _6798_ (.A1(net462),
    .A2(net1953),
    .A3(net312),
    .B1(_3550_),
    .X(_1061_));
 sky130_fd_sc_hd__and2_1 _6799_ (.A(net326),
    .B(net314),
    .X(_3551_));
 sky130_fd_sc_hd__a31o_1 _6800_ (.A1(net448),
    .A2(net1955),
    .A3(net313),
    .B1(_3551_),
    .X(_1062_));
 sky130_fd_sc_hd__and2_1 _6801_ (.A(net324),
    .B(net314),
    .X(_3552_));
 sky130_fd_sc_hd__a31o_1 _6802_ (.A1(net442),
    .A2(net1880),
    .A3(net313),
    .B1(_3552_),
    .X(_1063_));
 sky130_fd_sc_hd__and2_1 _6803_ (.A(net321),
    .B(net315),
    .X(_3553_));
 sky130_fd_sc_hd__a31o_1 _6804_ (.A1(net463),
    .A2(net1710),
    .A3(net312),
    .B1(_3553_),
    .X(_1064_));
 sky130_fd_sc_hd__and2_1 _6805_ (.A(net323),
    .B(net315),
    .X(_3554_));
 sky130_fd_sc_hd__a31o_1 _6806_ (.A1(net462),
    .A2(net1989),
    .A3(net312),
    .B1(_3554_),
    .X(_1065_));
 sky130_fd_sc_hd__and2_1 _6807_ (.A(net322),
    .B(net315),
    .X(_3555_));
 sky130_fd_sc_hd__a31o_1 _6808_ (.A1(net465),
    .A2(net1595),
    .A3(net312),
    .B1(_3555_),
    .X(_1066_));
 sky130_fd_sc_hd__and2_1 _6809_ (.A(net320),
    .B(net315),
    .X(_3556_));
 sky130_fd_sc_hd__a31o_1 _6810_ (.A1(net464),
    .A2(net1925),
    .A3(net312),
    .B1(_3556_),
    .X(_1067_));
 sky130_fd_sc_hd__and2_1 _6811_ (.A(net344),
    .B(net314),
    .X(_3557_));
 sky130_fd_sc_hd__a31o_1 _6812_ (.A1(net450),
    .A2(net1986),
    .A3(net313),
    .B1(_3557_),
    .X(_1068_));
 sky130_fd_sc_hd__nor2_1 _6813_ (.A(_1511_),
    .B(net312),
    .Y(_3558_));
 sky130_fd_sc_hd__a31o_1 _6814_ (.A1(net460),
    .A2(net1884),
    .A3(net312),
    .B1(_3558_),
    .X(_1069_));
 sky130_fd_sc_hd__and2_1 _6815_ (.A(net343),
    .B(net315),
    .X(_3559_));
 sky130_fd_sc_hd__a31o_1 _6816_ (.A1(net465),
    .A2(net1776),
    .A3(net312),
    .B1(_3559_),
    .X(_1070_));
 sky130_fd_sc_hd__and2_1 _6817_ (.A(net345),
    .B(net315),
    .X(_3560_));
 sky130_fd_sc_hd__a31o_1 _6818_ (.A1(net463),
    .A2(net1941),
    .A3(net312),
    .B1(_3560_),
    .X(_1071_));
 sky130_fd_sc_hd__and2_1 _6819_ (.A(net340),
    .B(net314),
    .X(_3561_));
 sky130_fd_sc_hd__a31o_1 _6820_ (.A1(net443),
    .A2(net1685),
    .A3(net313),
    .B1(_3561_),
    .X(_1072_));
 sky130_fd_sc_hd__and2_1 _6821_ (.A(net342),
    .B(net314),
    .X(_3562_));
 sky130_fd_sc_hd__a31o_1 _6822_ (.A1(net444),
    .A2(net1937),
    .A3(net313),
    .B1(_3562_),
    .X(_1073_));
 sky130_fd_sc_hd__and2_1 _6823_ (.A(net341),
    .B(net315),
    .X(_3563_));
 sky130_fd_sc_hd__a31o_1 _6824_ (.A1(net468),
    .A2(net1964),
    .A3(net312),
    .B1(_3563_),
    .X(_1074_));
 sky130_fd_sc_hd__and2_1 _6825_ (.A(net339),
    .B(net314),
    .X(_3564_));
 sky130_fd_sc_hd__a31o_1 _6826_ (.A1(net443),
    .A2(net1923),
    .A3(net313),
    .B1(_3564_),
    .X(_1075_));
 sky130_fd_sc_hd__and2_1 _6827_ (.A(net336),
    .B(net315),
    .X(_3565_));
 sky130_fd_sc_hd__a31o_1 _6828_ (.A1(net462),
    .A2(net1882),
    .A3(net312),
    .B1(_3565_),
    .X(_1076_));
 sky130_fd_sc_hd__and2_1 _6829_ (.A(net338),
    .B(net314),
    .X(_3566_));
 sky130_fd_sc_hd__a31o_1 _6830_ (.A1(net443),
    .A2(net1895),
    .A3(net313),
    .B1(_3566_),
    .X(_1077_));
 sky130_fd_sc_hd__and2_1 _6831_ (.A(net337),
    .B(net314),
    .X(_3567_));
 sky130_fd_sc_hd__a31o_1 _6832_ (.A1(net472),
    .A2(net1798),
    .A3(net313),
    .B1(_3567_),
    .X(_1078_));
 sky130_fd_sc_hd__and2_1 _6833_ (.A(net335),
    .B(net314),
    .X(_3568_));
 sky130_fd_sc_hd__a31o_1 _6834_ (.A1(net452),
    .A2(net1905),
    .A3(net313),
    .B1(_3568_),
    .X(_1079_));
 sky130_fd_sc_hd__and2_1 _6835_ (.A(net348),
    .B(net314),
    .X(_3569_));
 sky130_fd_sc_hd__a31o_1 _6836_ (.A1(net442),
    .A2(net1876),
    .A3(net313),
    .B1(_3569_),
    .X(_1080_));
 sky130_fd_sc_hd__and2_1 _6837_ (.A(net346),
    .B(net314),
    .X(_3570_));
 sky130_fd_sc_hd__a31o_1 _6838_ (.A1(net439),
    .A2(net1812),
    .A3(net313),
    .B1(_3570_),
    .X(_1081_));
 sky130_fd_sc_hd__and2_1 _6839_ (.A(net347),
    .B(net314),
    .X(_3571_));
 sky130_fd_sc_hd__a31o_1 _6840_ (.A1(net439),
    .A2(net1800),
    .A3(net313),
    .B1(_3571_),
    .X(_1082_));
 sky130_fd_sc_hd__and2_1 _6841_ (.A(net370),
    .B(net314),
    .X(_3572_));
 sky130_fd_sc_hd__a31o_1 _6842_ (.A1(net445),
    .A2(net1888),
    .A3(net313),
    .B1(_3572_),
    .X(_1083_));
 sky130_fd_sc_hd__nor2_4 _6843_ (.A(_2758_),
    .B(_3538_),
    .Y(_3573_));
 sky130_fd_sc_hd__or2_2 _6844_ (.A(_2758_),
    .B(_3538_),
    .X(_3574_));
 sky130_fd_sc_hd__nor2_2 _6845_ (.A(net479),
    .B(net257),
    .Y(_3575_));
 sky130_fd_sc_hd__nand2_1 _6846_ (.A(net470),
    .B(_3574_),
    .Y(_3576_));
 sky130_fd_sc_hd__o22a_1 _6847_ (.A1(net331),
    .A2(_3574_),
    .B1(_3576_),
    .B2(net980),
    .X(_1084_));
 sky130_fd_sc_hd__a22o_1 _6848_ (.A1(net332),
    .A2(net257),
    .B1(net220),
    .B2(net1443),
    .X(_1085_));
 sky130_fd_sc_hd__o22a_1 _6849_ (.A1(net333),
    .A2(_3574_),
    .B1(_3576_),
    .B2(net851),
    .X(_1086_));
 sky130_fd_sc_hd__a22o_1 _6850_ (.A1(net334),
    .A2(net257),
    .B1(net220),
    .B2(net1571),
    .X(_1087_));
 sky130_fd_sc_hd__a22o_1 _6851_ (.A1(net329),
    .A2(net257),
    .B1(net220),
    .B2(net1341),
    .X(_1088_));
 sky130_fd_sc_hd__a22o_1 _6852_ (.A1(_1741_),
    .A2(net257),
    .B1(net220),
    .B2(net1158),
    .X(_1089_));
 sky130_fd_sc_hd__a22o_1 _6853_ (.A1(net328),
    .A2(net257),
    .B1(net220),
    .B2(net1307),
    .X(_1090_));
 sky130_fd_sc_hd__a22o_1 _6854_ (.A1(net330),
    .A2(net256),
    .B1(net219),
    .B2(net1014),
    .X(_1091_));
 sky130_fd_sc_hd__a22o_1 _6855_ (.A1(net325),
    .A2(net256),
    .B1(net219),
    .B2(net1266),
    .X(_1092_));
 sky130_fd_sc_hd__a22o_1 _6856_ (.A1(net327),
    .A2(net257),
    .B1(net220),
    .B2(net1351),
    .X(_1093_));
 sky130_fd_sc_hd__a22o_1 _6857_ (.A1(net326),
    .A2(net256),
    .B1(net219),
    .B2(net1499),
    .X(_1094_));
 sky130_fd_sc_hd__a22o_1 _6858_ (.A1(net324),
    .A2(net256),
    .B1(net219),
    .B2(net1421),
    .X(_1095_));
 sky130_fd_sc_hd__a22o_1 _6859_ (.A1(_1821_),
    .A2(net257),
    .B1(net220),
    .B2(net1463),
    .X(_1096_));
 sky130_fd_sc_hd__a22o_1 _6860_ (.A1(net323),
    .A2(net257),
    .B1(net220),
    .B2(net1278),
    .X(_1097_));
 sky130_fd_sc_hd__a22o_1 _6861_ (.A1(net322),
    .A2(net257),
    .B1(net220),
    .B2(net1128),
    .X(_1098_));
 sky130_fd_sc_hd__a22o_1 _6862_ (.A1(net320),
    .A2(net257),
    .B1(net220),
    .B2(net936),
    .X(_1099_));
 sky130_fd_sc_hd__a22o_1 _6863_ (.A1(net344),
    .A2(net256),
    .B1(net219),
    .B2(net1605),
    .X(_1100_));
 sky130_fd_sc_hd__a22o_1 _6864_ (.A1(_1512_),
    .A2(net256),
    .B1(net219),
    .B2(net1699),
    .X(_1101_));
 sky130_fd_sc_hd__a22o_1 _6865_ (.A1(_1550_),
    .A2(net257),
    .B1(net220),
    .B2(net916),
    .X(_1102_));
 sky130_fd_sc_hd__a22o_1 _6866_ (.A1(net345),
    .A2(net257),
    .B1(net220),
    .B2(net1511),
    .X(_1103_));
 sky130_fd_sc_hd__a22o_1 _6867_ (.A1(net340),
    .A2(net256),
    .B1(net219),
    .B2(net958),
    .X(_1104_));
 sky130_fd_sc_hd__a22o_1 _6868_ (.A1(net342),
    .A2(net256),
    .B1(net219),
    .B2(net1473),
    .X(_1105_));
 sky130_fd_sc_hd__a22o_1 _6869_ (.A1(net341),
    .A2(net257),
    .B1(net220),
    .B2(net1469),
    .X(_1106_));
 sky130_fd_sc_hd__a22o_1 _6870_ (.A1(net339),
    .A2(net256),
    .B1(net219),
    .B2(net1172),
    .X(_1107_));
 sky130_fd_sc_hd__a22o_1 _6871_ (.A1(net336),
    .A2(net257),
    .B1(net220),
    .B2(net1585),
    .X(_1108_));
 sky130_fd_sc_hd__a22o_1 _6872_ (.A1(net338),
    .A2(net256),
    .B1(net219),
    .B2(net1311),
    .X(_1109_));
 sky130_fd_sc_hd__a22o_1 _6873_ (.A1(net337),
    .A2(net256),
    .B1(net219),
    .B2(net1427),
    .X(_1110_));
 sky130_fd_sc_hd__a22o_1 _6874_ (.A1(net335),
    .A2(net256),
    .B1(net219),
    .B2(net1419),
    .X(_1111_));
 sky130_fd_sc_hd__a22o_1 _6875_ (.A1(_1473_),
    .A2(net256),
    .B1(net219),
    .B2(net1758),
    .X(_1112_));
 sky130_fd_sc_hd__a22o_1 _6876_ (.A1(net346),
    .A2(net256),
    .B1(net219),
    .B2(net1483),
    .X(_1113_));
 sky130_fd_sc_hd__a22o_1 _6877_ (.A1(net347),
    .A2(net256),
    .B1(net219),
    .B2(net1465),
    .X(_1114_));
 sky130_fd_sc_hd__a22o_1 _6878_ (.A1(net370),
    .A2(net256),
    .B1(net219),
    .B2(net1268),
    .X(_1115_));
 sky130_fd_sc_hd__or2_2 _6879_ (.A(net365),
    .B(_2753_),
    .X(_3577_));
 sky130_fd_sc_hd__nor2_4 _6880_ (.A(_2767_),
    .B(_3577_),
    .Y(_3578_));
 sky130_fd_sc_hd__or2_1 _6881_ (.A(_2767_),
    .B(_3577_),
    .X(_3579_));
 sky130_fd_sc_hd__nor2_4 _6882_ (.A(net473),
    .B(net254),
    .Y(_3580_));
 sky130_fd_sc_hd__nand2_1 _6883_ (.A(net467),
    .B(_3579_),
    .Y(_3581_));
 sky130_fd_sc_hd__o22a_1 _6884_ (.A1(net331),
    .A2(_3579_),
    .B1(_3581_),
    .B2(net890),
    .X(_1116_));
 sky130_fd_sc_hd__o22a_1 _6885_ (.A1(net332),
    .A2(_3579_),
    .B1(_3581_),
    .B2(net876),
    .X(_1117_));
 sky130_fd_sc_hd__a22o_1 _6886_ (.A1(net333),
    .A2(net255),
    .B1(net218),
    .B2(net1052),
    .X(_1118_));
 sky130_fd_sc_hd__o22a_1 _6887_ (.A1(net334),
    .A2(_3579_),
    .B1(_3581_),
    .B2(net878),
    .X(_1119_));
 sky130_fd_sc_hd__a22o_1 _6888_ (.A1(net329),
    .A2(net255),
    .B1(net218),
    .B2(net1569),
    .X(_1120_));
 sky130_fd_sc_hd__a22o_1 _6889_ (.A1(_1741_),
    .A2(net255),
    .B1(net218),
    .B2(net1200),
    .X(_1121_));
 sky130_fd_sc_hd__a22o_1 _6890_ (.A1(net328),
    .A2(net255),
    .B1(net218),
    .B2(net1505),
    .X(_1122_));
 sky130_fd_sc_hd__a22o_1 _6891_ (.A1(net330),
    .A2(net254),
    .B1(net217),
    .B2(net1234),
    .X(_1123_));
 sky130_fd_sc_hd__a22o_1 _6892_ (.A1(net325),
    .A2(net254),
    .B1(net217),
    .B2(net1050),
    .X(_1124_));
 sky130_fd_sc_hd__a22o_1 _6893_ (.A1(net327),
    .A2(net255),
    .B1(net218),
    .B2(net1481),
    .X(_1125_));
 sky130_fd_sc_hd__a22o_1 _6894_ (.A1(net326),
    .A2(net254),
    .B1(net217),
    .B2(net1222),
    .X(_1126_));
 sky130_fd_sc_hd__a22o_1 _6895_ (.A1(net324),
    .A2(net254),
    .B1(net217),
    .B2(net1317),
    .X(_1127_));
 sky130_fd_sc_hd__a22o_1 _6896_ (.A1(net321),
    .A2(net255),
    .B1(net218),
    .B2(net1068),
    .X(_1128_));
 sky130_fd_sc_hd__a22o_1 _6897_ (.A1(_1800_),
    .A2(net255),
    .B1(net218),
    .B2(net1323),
    .X(_1129_));
 sky130_fd_sc_hd__a22o_1 _6898_ (.A1(net322),
    .A2(net255),
    .B1(net218),
    .B2(net1284),
    .X(_1130_));
 sky130_fd_sc_hd__a22o_1 _6899_ (.A1(net320),
    .A2(net255),
    .B1(net218),
    .B2(net1517),
    .X(_1131_));
 sky130_fd_sc_hd__a22o_1 _6900_ (.A1(net344),
    .A2(net254),
    .B1(net217),
    .B2(net1335),
    .X(_1132_));
 sky130_fd_sc_hd__a22o_1 _6901_ (.A1(_1512_),
    .A2(net255),
    .B1(net217),
    .B2(net1122),
    .X(_1133_));
 sky130_fd_sc_hd__a22o_1 _6902_ (.A1(net343),
    .A2(net255),
    .B1(net218),
    .B2(net1178),
    .X(_1134_));
 sky130_fd_sc_hd__a22o_1 _6903_ (.A1(net345),
    .A2(net255),
    .B1(net218),
    .B2(net1002),
    .X(_1135_));
 sky130_fd_sc_hd__a22o_1 _6904_ (.A1(net340),
    .A2(net254),
    .B1(net217),
    .B2(net1523),
    .X(_1136_));
 sky130_fd_sc_hd__a22o_1 _6905_ (.A1(net342),
    .A2(net254),
    .B1(net217),
    .B2(net1449),
    .X(_1137_));
 sky130_fd_sc_hd__a22o_1 _6906_ (.A1(net341),
    .A2(net255),
    .B1(net218),
    .B2(net1535),
    .X(_1138_));
 sky130_fd_sc_hd__a22o_1 _6907_ (.A1(net339),
    .A2(net254),
    .B1(net217),
    .B2(net1701),
    .X(_1139_));
 sky130_fd_sc_hd__a22o_1 _6908_ (.A1(net336),
    .A2(net255),
    .B1(net218),
    .B2(net1118),
    .X(_1140_));
 sky130_fd_sc_hd__a22o_1 _6909_ (.A1(net338),
    .A2(net254),
    .B1(net217),
    .B2(net1299),
    .X(_1141_));
 sky130_fd_sc_hd__a22o_1 _6910_ (.A1(net337),
    .A2(net254),
    .B1(net217),
    .B2(net1054),
    .X(_1142_));
 sky130_fd_sc_hd__a22o_1 _6911_ (.A1(net335),
    .A2(net254),
    .B1(net217),
    .B2(net1290),
    .X(_1143_));
 sky130_fd_sc_hd__a22o_1 _6912_ (.A1(net348),
    .A2(net254),
    .B1(net217),
    .B2(net1423),
    .X(_1144_));
 sky130_fd_sc_hd__a22o_1 _6913_ (.A1(net346),
    .A2(net254),
    .B1(net217),
    .B2(net1381),
    .X(_1145_));
 sky130_fd_sc_hd__a22o_1 _6914_ (.A1(net347),
    .A2(net254),
    .B1(net217),
    .B2(net1718),
    .X(_1146_));
 sky130_fd_sc_hd__a22o_1 _6915_ (.A1(net370),
    .A2(net254),
    .B1(net217),
    .B2(net1788),
    .X(_1147_));
 sky130_fd_sc_hd__nor2_2 _6916_ (.A(_2743_),
    .B(_3577_),
    .Y(_3582_));
 sky130_fd_sc_hd__or2_4 _6917_ (.A(_2743_),
    .B(_3577_),
    .X(_3583_));
 sky130_fd_sc_hd__and2_1 _6918_ (.A(net331),
    .B(net253),
    .X(_3584_));
 sky130_fd_sc_hd__a31o_1 _6919_ (.A1(net468),
    .A2(net1786),
    .A3(net250),
    .B1(_3584_),
    .X(_1148_));
 sky130_fd_sc_hd__and2_1 _6920_ (.A(net332),
    .B(net253),
    .X(_3585_));
 sky130_fd_sc_hd__a31o_1 _6921_ (.A1(net467),
    .A2(net1774),
    .A3(net250),
    .B1(_3585_),
    .X(_1149_));
 sky130_fd_sc_hd__and2_1 _6922_ (.A(net333),
    .B(net253),
    .X(_3586_));
 sky130_fd_sc_hd__a31o_1 _6923_ (.A1(net468),
    .A2(net1826),
    .A3(net250),
    .B1(_3586_),
    .X(_1150_));
 sky130_fd_sc_hd__or3_1 _6924_ (.A(net481),
    .B(net2129),
    .C(net253),
    .X(_3587_));
 sky130_fd_sc_hd__o21a_1 _6925_ (.A1(net334),
    .A2(net250),
    .B1(_3587_),
    .X(_1151_));
 sky130_fd_sc_hd__and2_1 _6926_ (.A(net329),
    .B(net252),
    .X(_3588_));
 sky130_fd_sc_hd__a31o_1 _6927_ (.A1(net463),
    .A2(net1838),
    .A3(net250),
    .B1(_3588_),
    .X(_1152_));
 sky130_fd_sc_hd__nor2_1 _6928_ (.A(_1740_),
    .B(_3583_),
    .Y(_3589_));
 sky130_fd_sc_hd__a31o_1 _6929_ (.A1(net464),
    .A2(net1897),
    .A3(_3583_),
    .B1(_3589_),
    .X(_1153_));
 sky130_fd_sc_hd__and2_1 _6930_ (.A(net328),
    .B(net252),
    .X(_3590_));
 sky130_fd_sc_hd__a31o_1 _6931_ (.A1(net460),
    .A2(net1931),
    .A3(net250),
    .B1(_3590_),
    .X(_1154_));
 sky130_fd_sc_hd__and2_1 _6932_ (.A(net330),
    .B(net252),
    .X(_3591_));
 sky130_fd_sc_hd__a31o_1 _6933_ (.A1(net439),
    .A2(net1886),
    .A3(net251),
    .B1(_3591_),
    .X(_1155_));
 sky130_fd_sc_hd__and2_1 _6934_ (.A(net325),
    .B(net252),
    .X(_3592_));
 sky130_fd_sc_hd__a31o_1 _6935_ (.A1(net441),
    .A2(net1742),
    .A3(net251),
    .B1(_3592_),
    .X(_1156_));
 sky130_fd_sc_hd__and2_1 _6936_ (.A(net327),
    .B(net253),
    .X(_3593_));
 sky130_fd_sc_hd__a31o_1 _6937_ (.A1(net462),
    .A2(net1911),
    .A3(net250),
    .B1(_3593_),
    .X(_1157_));
 sky130_fd_sc_hd__and2_1 _6938_ (.A(net326),
    .B(net252),
    .X(_3594_));
 sky130_fd_sc_hd__a31o_1 _6939_ (.A1(net448),
    .A2(net1655),
    .A3(net251),
    .B1(_3594_),
    .X(_1158_));
 sky130_fd_sc_hd__and2_1 _6940_ (.A(net324),
    .B(net252),
    .X(_3595_));
 sky130_fd_sc_hd__a31o_1 _6941_ (.A1(net442),
    .A2(net1617),
    .A3(net251),
    .B1(_3595_),
    .X(_1159_));
 sky130_fd_sc_hd__and2_1 _6942_ (.A(net321),
    .B(net253),
    .X(_3596_));
 sky130_fd_sc_hd__a31o_1 _6943_ (.A1(net463),
    .A2(net1913),
    .A3(net250),
    .B1(_3596_),
    .X(_1160_));
 sky130_fd_sc_hd__and2_1 _6944_ (.A(net323),
    .B(net253),
    .X(_3597_));
 sky130_fd_sc_hd__a31o_1 _6945_ (.A1(net463),
    .A2(net1907),
    .A3(net250),
    .B1(_3597_),
    .X(_1161_));
 sky130_fd_sc_hd__and2_1 _6946_ (.A(net322),
    .B(net253),
    .X(_3598_));
 sky130_fd_sc_hd__a31o_1 _6947_ (.A1(net464),
    .A2(net1959),
    .A3(net250),
    .B1(_3598_),
    .X(_1162_));
 sky130_fd_sc_hd__and2_1 _6948_ (.A(net320),
    .B(net253),
    .X(_3599_));
 sky130_fd_sc_hd__a31o_1 _6949_ (.A1(net458),
    .A2(net1659),
    .A3(net250),
    .B1(_3599_),
    .X(_1163_));
 sky130_fd_sc_hd__and2_1 _6950_ (.A(net344),
    .B(net252),
    .X(_3600_));
 sky130_fd_sc_hd__a31o_1 _6951_ (.A1(net452),
    .A2(net1978),
    .A3(net251),
    .B1(_3600_),
    .X(_1164_));
 sky130_fd_sc_hd__nor2_1 _6952_ (.A(_1511_),
    .B(net250),
    .Y(_3601_));
 sky130_fd_sc_hd__a31o_1 _6953_ (.A1(net460),
    .A2(net1961),
    .A3(net250),
    .B1(_3601_),
    .X(_1165_));
 sky130_fd_sc_hd__and2_1 _6954_ (.A(net343),
    .B(net253),
    .X(_3602_));
 sky130_fd_sc_hd__a31o_1 _6955_ (.A1(net471),
    .A2(net1929),
    .A3(net250),
    .B1(_3602_),
    .X(_1166_));
 sky130_fd_sc_hd__and2_1 _6956_ (.A(_1526_),
    .B(net253),
    .X(_3603_));
 sky130_fd_sc_hd__a31o_1 _6957_ (.A1(net467),
    .A2(net1943),
    .A3(net250),
    .B1(_3603_),
    .X(_1167_));
 sky130_fd_sc_hd__and2_1 _6958_ (.A(net340),
    .B(net252),
    .X(_3604_));
 sky130_fd_sc_hd__a31o_1 _6959_ (.A1(net444),
    .A2(net1639),
    .A3(net251),
    .B1(_3604_),
    .X(_1168_));
 sky130_fd_sc_hd__and2_1 _6960_ (.A(net342),
    .B(net252),
    .X(_3605_));
 sky130_fd_sc_hd__a31o_1 _6961_ (.A1(net444),
    .A2(net1770),
    .A3(net251),
    .B1(_3605_),
    .X(_1169_));
 sky130_fd_sc_hd__and2_1 _6962_ (.A(net341),
    .B(net253),
    .X(_3606_));
 sky130_fd_sc_hd__a31o_1 _6963_ (.A1(net468),
    .A2(net1966),
    .A3(net251),
    .B1(_3606_),
    .X(_1170_));
 sky130_fd_sc_hd__and2_1 _6964_ (.A(net339),
    .B(net252),
    .X(_3607_));
 sky130_fd_sc_hd__a31o_1 _6965_ (.A1(net443),
    .A2(net1844),
    .A3(net251),
    .B1(_3607_),
    .X(_1171_));
 sky130_fd_sc_hd__and2_1 _6966_ (.A(net336),
    .B(net253),
    .X(_3608_));
 sky130_fd_sc_hd__a31o_1 _6967_ (.A1(net463),
    .A2(net1976),
    .A3(_3583_),
    .B1(_3608_),
    .X(_1172_));
 sky130_fd_sc_hd__and2_1 _6968_ (.A(net338),
    .B(net252),
    .X(_3609_));
 sky130_fd_sc_hd__a31o_1 _6969_ (.A1(net443),
    .A2(net1868),
    .A3(net251),
    .B1(_3609_),
    .X(_1173_));
 sky130_fd_sc_hd__and2_1 _6970_ (.A(net337),
    .B(net252),
    .X(_3610_));
 sky130_fd_sc_hd__a31o_1 _6971_ (.A1(net443),
    .A2(net1927),
    .A3(net251),
    .B1(_3610_),
    .X(_1174_));
 sky130_fd_sc_hd__and2_1 _6972_ (.A(net335),
    .B(net253),
    .X(_3611_));
 sky130_fd_sc_hd__a31o_1 _6973_ (.A1(net452),
    .A2(net1980),
    .A3(net250),
    .B1(_3611_),
    .X(_1175_));
 sky130_fd_sc_hd__and2_1 _6974_ (.A(net348),
    .B(net252),
    .X(_3612_));
 sky130_fd_sc_hd__a31o_1 _6975_ (.A1(net439),
    .A2(net1903),
    .A3(net251),
    .B1(_3612_),
    .X(_1176_));
 sky130_fd_sc_hd__and2_1 _6976_ (.A(net346),
    .B(net252),
    .X(_3613_));
 sky130_fd_sc_hd__a31o_1 _6977_ (.A1(net439),
    .A2(net1808),
    .A3(net251),
    .B1(_3613_),
    .X(_1177_));
 sky130_fd_sc_hd__and2_1 _6978_ (.A(net347),
    .B(net252),
    .X(_3614_));
 sky130_fd_sc_hd__a31o_1 _6979_ (.A1(net439),
    .A2(net1957),
    .A3(net251),
    .B1(_3614_),
    .X(_1178_));
 sky130_fd_sc_hd__and2_1 _6980_ (.A(net370),
    .B(net252),
    .X(_3615_));
 sky130_fd_sc_hd__a31o_1 _6981_ (.A1(net445),
    .A2(net1862),
    .A3(net251),
    .B1(_3615_),
    .X(_1179_));
 sky130_fd_sc_hd__nor3_4 _6982_ (.A(net365),
    .B(_2767_),
    .C(_3538_),
    .Y(_3616_));
 sky130_fd_sc_hd__or3_2 _6983_ (.A(_2744_),
    .B(_2767_),
    .C(_3538_),
    .X(_3617_));
 sky130_fd_sc_hd__nor2_4 _6984_ (.A(net473),
    .B(net310),
    .Y(_3618_));
 sky130_fd_sc_hd__nand2_1 _6985_ (.A(net471),
    .B(_3617_),
    .Y(_3619_));
 sky130_fd_sc_hd__o22a_1 _6986_ (.A1(net331),
    .A2(_3617_),
    .B1(_3619_),
    .B2(net910),
    .X(_1180_));
 sky130_fd_sc_hd__o22a_1 _6987_ (.A1(net332),
    .A2(_3617_),
    .B1(_3619_),
    .B2(net864),
    .X(_1181_));
 sky130_fd_sc_hd__o22a_1 _6988_ (.A1(net333),
    .A2(_3617_),
    .B1(_3619_),
    .B2(net888),
    .X(_1182_));
 sky130_fd_sc_hd__a22o_1 _6989_ (.A1(net334),
    .A2(net311),
    .B1(net249),
    .B2(net1379),
    .X(_1183_));
 sky130_fd_sc_hd__a22o_1 _6990_ (.A1(net329),
    .A2(net311),
    .B1(net249),
    .B2(net1212),
    .X(_1184_));
 sky130_fd_sc_hd__a22o_1 _6991_ (.A1(_1741_),
    .A2(net311),
    .B1(net249),
    .B2(net1274),
    .X(_1185_));
 sky130_fd_sc_hd__a22o_1 _6992_ (.A1(net328),
    .A2(net311),
    .B1(net249),
    .B2(net1162),
    .X(_1186_));
 sky130_fd_sc_hd__a22o_1 _6993_ (.A1(net330),
    .A2(net310),
    .B1(net248),
    .B2(net1282),
    .X(_1187_));
 sky130_fd_sc_hd__a22o_1 _6994_ (.A1(net325),
    .A2(net310),
    .B1(net248),
    .B2(net1467),
    .X(_1188_));
 sky130_fd_sc_hd__a22o_1 _6995_ (.A1(net327),
    .A2(net311),
    .B1(net249),
    .B2(net1116),
    .X(_1189_));
 sky130_fd_sc_hd__a22o_1 _6996_ (.A1(net326),
    .A2(net310),
    .B1(net248),
    .B2(net1583),
    .X(_1190_));
 sky130_fd_sc_hd__a22o_1 _6997_ (.A1(net324),
    .A2(net310),
    .B1(net248),
    .B2(net1475),
    .X(_1191_));
 sky130_fd_sc_hd__a22o_1 _6998_ (.A1(net321),
    .A2(net311),
    .B1(net249),
    .B2(net1100),
    .X(_1192_));
 sky130_fd_sc_hd__a22o_1 _6999_ (.A1(net323),
    .A2(net311),
    .B1(net249),
    .B2(net1802),
    .X(_1193_));
 sky130_fd_sc_hd__a22o_1 _7000_ (.A1(net322),
    .A2(net311),
    .B1(net249),
    .B2(net972),
    .X(_1194_));
 sky130_fd_sc_hd__a22o_1 _7001_ (.A1(net320),
    .A2(net311),
    .B1(net249),
    .B2(net1521),
    .X(_1195_));
 sky130_fd_sc_hd__a22o_1 _7002_ (.A1(net344),
    .A2(net310),
    .B1(net248),
    .B2(net1373),
    .X(_1196_));
 sky130_fd_sc_hd__a22o_1 _7003_ (.A1(_1512_),
    .A2(net311),
    .B1(net248),
    .B2(net1345),
    .X(_1197_));
 sky130_fd_sc_hd__a22o_1 _7004_ (.A1(net343),
    .A2(net311),
    .B1(net249),
    .B2(net1088),
    .X(_1198_));
 sky130_fd_sc_hd__a22o_1 _7005_ (.A1(net345),
    .A2(net311),
    .B1(net249),
    .B2(net1355),
    .X(_1199_));
 sky130_fd_sc_hd__a22o_1 _7006_ (.A1(net340),
    .A2(net310),
    .B1(net248),
    .B2(net1295),
    .X(_1200_));
 sky130_fd_sc_hd__a22o_1 _7007_ (.A1(net342),
    .A2(net310),
    .B1(net248),
    .B2(net1383),
    .X(_1201_));
 sky130_fd_sc_hd__a22o_1 _7008_ (.A1(net341),
    .A2(net311),
    .B1(net249),
    .B2(net1790),
    .X(_1202_));
 sky130_fd_sc_hd__a22o_1 _7009_ (.A1(net339),
    .A2(net310),
    .B1(net248),
    .B2(net1417),
    .X(_1203_));
 sky130_fd_sc_hd__a22o_1 _7010_ (.A1(net336),
    .A2(net311),
    .B1(net249),
    .B2(net1272),
    .X(_1204_));
 sky130_fd_sc_hd__a22o_1 _7011_ (.A1(net338),
    .A2(net310),
    .B1(net248),
    .B2(net1126),
    .X(_1205_));
 sky130_fd_sc_hd__a22o_1 _7012_ (.A1(net337),
    .A2(net310),
    .B1(net248),
    .B2(net1012),
    .X(_1206_));
 sky130_fd_sc_hd__a22o_1 _7013_ (.A1(net335),
    .A2(net310),
    .B1(net248),
    .B2(net1730),
    .X(_1207_));
 sky130_fd_sc_hd__a22o_1 _7014_ (.A1(net348),
    .A2(net310),
    .B1(net248),
    .B2(net998),
    .X(_1208_));
 sky130_fd_sc_hd__a22o_1 _7015_ (.A1(net346),
    .A2(net310),
    .B1(net248),
    .B2(net1567),
    .X(_1209_));
 sky130_fd_sc_hd__a22o_1 _7016_ (.A1(net347),
    .A2(net310),
    .B1(net248),
    .B2(net898),
    .X(_1210_));
 sky130_fd_sc_hd__a22o_1 _7017_ (.A1(net370),
    .A2(net310),
    .B1(net248),
    .B2(net1321),
    .X(_1211_));
 sky130_fd_sc_hd__nor2_4 _7018_ (.A(_2752_),
    .B(_3538_),
    .Y(_3620_));
 sky130_fd_sc_hd__or2_1 _7019_ (.A(_2752_),
    .B(_3538_),
    .X(_3621_));
 sky130_fd_sc_hd__nor2_4 _7020_ (.A(net473),
    .B(net246),
    .Y(_3622_));
 sky130_fd_sc_hd__nand2_1 _7021_ (.A(net470),
    .B(_3621_),
    .Y(_3623_));
 sky130_fd_sc_hd__a22o_1 _7022_ (.A1(net331),
    .A2(net247),
    .B1(net216),
    .B2(net1016),
    .X(_1212_));
 sky130_fd_sc_hd__o22a_1 _7023_ (.A1(net332),
    .A2(_3621_),
    .B1(_3623_),
    .B2(net1010),
    .X(_1213_));
 sky130_fd_sc_hd__o22a_1 _7024_ (.A1(net333),
    .A2(_3621_),
    .B1(_3623_),
    .B2(net950),
    .X(_1214_));
 sky130_fd_sc_hd__a22o_1 _7025_ (.A1(net334),
    .A2(net247),
    .B1(net216),
    .B2(net1411),
    .X(_1215_));
 sky130_fd_sc_hd__a22o_1 _7026_ (.A1(net329),
    .A2(net247),
    .B1(net216),
    .B2(net938),
    .X(_1216_));
 sky130_fd_sc_hd__a22o_1 _7027_ (.A1(_1741_),
    .A2(net247),
    .B1(net216),
    .B2(net1407),
    .X(_1217_));
 sky130_fd_sc_hd__a22o_1 _7028_ (.A1(net328),
    .A2(net247),
    .B1(net216),
    .B2(net1471),
    .X(_1218_));
 sky130_fd_sc_hd__a22o_1 _7029_ (.A1(net330),
    .A2(net246),
    .B1(net215),
    .B2(net1146),
    .X(_1219_));
 sky130_fd_sc_hd__a22o_1 _7030_ (.A1(net325),
    .A2(net246),
    .B1(net215),
    .B2(net1613),
    .X(_1220_));
 sky130_fd_sc_hd__a22o_1 _7031_ (.A1(net327),
    .A2(net247),
    .B1(net216),
    .B2(net1192),
    .X(_1221_));
 sky130_fd_sc_hd__a22o_1 _7032_ (.A1(net326),
    .A2(net246),
    .B1(net215),
    .B2(net1609),
    .X(_1222_));
 sky130_fd_sc_hd__a22o_1 _7033_ (.A1(net324),
    .A2(net246),
    .B1(net215),
    .B2(net1112),
    .X(_1223_));
 sky130_fd_sc_hd__a22o_1 _7034_ (.A1(net321),
    .A2(net247),
    .B1(net216),
    .B2(net1018),
    .X(_1224_));
 sky130_fd_sc_hd__a22o_1 _7035_ (.A1(net323),
    .A2(net247),
    .B1(net216),
    .B2(net1661),
    .X(_1225_));
 sky130_fd_sc_hd__a22o_1 _7036_ (.A1(net322),
    .A2(net247),
    .B1(net216),
    .B2(net954),
    .X(_1226_));
 sky130_fd_sc_hd__a22o_1 _7037_ (.A1(net320),
    .A2(net247),
    .B1(net216),
    .B2(net1705),
    .X(_1227_));
 sky130_fd_sc_hd__a22o_1 _7038_ (.A1(net344),
    .A2(net246),
    .B1(net215),
    .B2(net1543),
    .X(_1228_));
 sky130_fd_sc_hd__a22o_1 _7039_ (.A1(_1512_),
    .A2(net247),
    .B1(net215),
    .B2(net1092),
    .X(_1229_));
 sky130_fd_sc_hd__a22o_1 _7040_ (.A1(net343),
    .A2(net247),
    .B1(net216),
    .B2(net1363),
    .X(_1230_));
 sky130_fd_sc_hd__a22o_1 _7041_ (.A1(net345),
    .A2(net247),
    .B1(net216),
    .B2(net1738),
    .X(_1231_));
 sky130_fd_sc_hd__a22o_1 _7042_ (.A1(net340),
    .A2(net246),
    .B1(net215),
    .B2(net1371),
    .X(_1232_));
 sky130_fd_sc_hd__a22o_1 _7043_ (.A1(net342),
    .A2(net246),
    .B1(net215),
    .B2(net1006),
    .X(_1233_));
 sky130_fd_sc_hd__a22o_1 _7044_ (.A1(net341),
    .A2(net247),
    .B1(net216),
    .B2(net1445),
    .X(_1234_));
 sky130_fd_sc_hd__a22o_1 _7045_ (.A1(net339),
    .A2(net246),
    .B1(net215),
    .B2(net1286),
    .X(_1235_));
 sky130_fd_sc_hd__a22o_1 _7046_ (.A1(net336),
    .A2(net247),
    .B1(net216),
    .B2(net1226),
    .X(_1236_));
 sky130_fd_sc_hd__a22o_1 _7047_ (.A1(net338),
    .A2(net246),
    .B1(net215),
    .B2(net1365),
    .X(_1237_));
 sky130_fd_sc_hd__a22o_1 _7048_ (.A1(net337),
    .A2(net246),
    .B1(net215),
    .B2(net994),
    .X(_1238_));
 sky130_fd_sc_hd__a22o_1 _7049_ (.A1(net335),
    .A2(net246),
    .B1(net215),
    .B2(net1581),
    .X(_1239_));
 sky130_fd_sc_hd__a22o_1 _7050_ (.A1(net348),
    .A2(net246),
    .B1(net215),
    .B2(net1136),
    .X(_1240_));
 sky130_fd_sc_hd__a22o_1 _7051_ (.A1(net346),
    .A2(net246),
    .B1(net215),
    .B2(net1764),
    .X(_1241_));
 sky130_fd_sc_hd__a22o_1 _7052_ (.A1(net347),
    .A2(net246),
    .B1(net215),
    .B2(net966),
    .X(_1242_));
 sky130_fd_sc_hd__a22o_1 _7053_ (.A1(net370),
    .A2(net246),
    .B1(net215),
    .B2(net1240),
    .X(_1243_));
 sky130_fd_sc_hd__nor3_1 _7054_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2752_),
    .Y(_3624_));
 sky130_fd_sc_hd__or3_4 _7055_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2752_),
    .X(_3625_));
 sky130_fd_sc_hd__and2_1 _7056_ (.A(net331),
    .B(net245),
    .X(_3626_));
 sky130_fd_sc_hd__a31o_1 _7057_ (.A1(net468),
    .A2(net1760),
    .A3(net242),
    .B1(_3626_),
    .X(_1274_));
 sky130_fd_sc_hd__or3_1 _7058_ (.A(net481),
    .B(net2114),
    .C(net244),
    .X(_3627_));
 sky130_fd_sc_hd__o21a_1 _7059_ (.A1(net332),
    .A2(net242),
    .B1(_3627_),
    .X(_1275_));
 sky130_fd_sc_hd__and2_1 _7060_ (.A(net333),
    .B(net244),
    .X(_3628_));
 sky130_fd_sc_hd__a31o_1 _7061_ (.A1(net470),
    .A2(net1878),
    .A3(_3625_),
    .B1(_3628_),
    .X(_1276_));
 sky130_fd_sc_hd__and2_1 _7062_ (.A(net334),
    .B(net244),
    .X(_3629_));
 sky130_fd_sc_hd__a31o_1 _7063_ (.A1(net470),
    .A2(net1852),
    .A3(net242),
    .B1(_3629_),
    .X(_1277_));
 sky130_fd_sc_hd__and2_1 _7064_ (.A(net329),
    .B(net244),
    .X(_3630_));
 sky130_fd_sc_hd__a31o_1 _7065_ (.A1(net463),
    .A2(net1933),
    .A3(_3625_),
    .B1(_3630_),
    .X(_1278_));
 sky130_fd_sc_hd__or3b_1 _7066_ (.A(net480),
    .B(net244),
    .C_N(net2148),
    .X(_3631_));
 sky130_fd_sc_hd__o21ai_1 _7067_ (.A1(_1740_),
    .A2(net242),
    .B1(_3631_),
    .Y(_1279_));
 sky130_fd_sc_hd__and2_1 _7068_ (.A(net328),
    .B(net244),
    .X(_3632_));
 sky130_fd_sc_hd__a31o_1 _7069_ (.A1(net460),
    .A2(net1848),
    .A3(net242),
    .B1(_3632_),
    .X(_1280_));
 sky130_fd_sc_hd__and2_1 _7070_ (.A(net330),
    .B(net245),
    .X(_3633_));
 sky130_fd_sc_hd__a31o_1 _7071_ (.A1(net440),
    .A2(net1856),
    .A3(net243),
    .B1(_3633_),
    .X(_1281_));
 sky130_fd_sc_hd__and2_1 _7072_ (.A(net325),
    .B(net245),
    .X(_3634_));
 sky130_fd_sc_hd__a31o_1 _7073_ (.A1(net447),
    .A2(net1970),
    .A3(net243),
    .B1(_3634_),
    .X(_1282_));
 sky130_fd_sc_hd__and2_1 _7074_ (.A(net327),
    .B(net244),
    .X(_3635_));
 sky130_fd_sc_hd__a31o_1 _7075_ (.A1(net460),
    .A2(net1754),
    .A3(net242),
    .B1(_3635_),
    .X(_1283_));
 sky130_fd_sc_hd__and2_1 _7076_ (.A(_1767_),
    .B(net245),
    .X(_3636_));
 sky130_fd_sc_hd__a31o_1 _7077_ (.A1(net449),
    .A2(net1840),
    .A3(net243),
    .B1(_3636_),
    .X(_1284_));
 sky130_fd_sc_hd__and2_1 _7078_ (.A(net324),
    .B(net245),
    .X(_3637_));
 sky130_fd_sc_hd__a31o_1 _7079_ (.A1(net441),
    .A2(net1951),
    .A3(net243),
    .B1(_3637_),
    .X(_1285_));
 sky130_fd_sc_hd__and2_1 _7080_ (.A(net321),
    .B(net244),
    .X(_3638_));
 sky130_fd_sc_hd__a31o_1 _7081_ (.A1(net463),
    .A2(net1667),
    .A3(net242),
    .B1(_3638_),
    .X(_1286_));
 sky130_fd_sc_hd__and2_1 _7082_ (.A(net323),
    .B(net244),
    .X(_3639_));
 sky130_fd_sc_hd__a31o_1 _7083_ (.A1(net462),
    .A2(net1994),
    .A3(net242),
    .B1(_3639_),
    .X(_1287_));
 sky130_fd_sc_hd__and2_1 _7084_ (.A(net322),
    .B(net244),
    .X(_3640_));
 sky130_fd_sc_hd__a31o_1 _7085_ (.A1(net471),
    .A2(net1909),
    .A3(net242),
    .B1(_3640_),
    .X(_1288_));
 sky130_fd_sc_hd__and2_1 _7086_ (.A(net320),
    .B(net244),
    .X(_3641_));
 sky130_fd_sc_hd__a31o_1 _7087_ (.A1(net457),
    .A2(net1814),
    .A3(net242),
    .B1(_3641_),
    .X(_1289_));
 sky130_fd_sc_hd__and2_1 _7088_ (.A(net344),
    .B(net245),
    .X(_3642_));
 sky130_fd_sc_hd__a31o_1 _7089_ (.A1(net452),
    .A2(net1935),
    .A3(net243),
    .B1(_3642_),
    .X(_1290_));
 sky130_fd_sc_hd__nor2_1 _7090_ (.A(_1511_),
    .B(net242),
    .Y(_3643_));
 sky130_fd_sc_hd__a31o_1 _7091_ (.A1(net452),
    .A2(net1671),
    .A3(net243),
    .B1(_3643_),
    .X(_1291_));
 sky130_fd_sc_hd__and2_1 _7092_ (.A(net343),
    .B(net244),
    .X(_3644_));
 sky130_fd_sc_hd__a31o_1 _7093_ (.A1(net465),
    .A2(net1714),
    .A3(net242),
    .B1(_3644_),
    .X(_1292_));
 sky130_fd_sc_hd__and2_1 _7094_ (.A(net345),
    .B(net244),
    .X(_3645_));
 sky130_fd_sc_hd__a31o_1 _7095_ (.A1(net464),
    .A2(net1870),
    .A3(net242),
    .B1(_3645_),
    .X(_1293_));
 sky130_fd_sc_hd__and2_1 _7096_ (.A(net340),
    .B(net245),
    .X(_3646_));
 sky130_fd_sc_hd__a31o_1 _7097_ (.A1(net443),
    .A2(net1820),
    .A3(net243),
    .B1(_3646_),
    .X(_1294_));
 sky130_fd_sc_hd__and2_1 _7098_ (.A(net342),
    .B(net245),
    .X(_3647_));
 sky130_fd_sc_hd__a31o_1 _7099_ (.A1(net444),
    .A2(net1866),
    .A3(net243),
    .B1(_3647_),
    .X(_1295_));
 sky130_fd_sc_hd__and2_1 _7100_ (.A(net341),
    .B(net244),
    .X(_3648_));
 sky130_fd_sc_hd__a31o_1 _7101_ (.A1(net467),
    .A2(net1832),
    .A3(net242),
    .B1(_3648_),
    .X(_1296_));
 sky130_fd_sc_hd__and2_1 _7102_ (.A(net339),
    .B(net245),
    .X(_3649_));
 sky130_fd_sc_hd__a31o_1 _7103_ (.A1(net443),
    .A2(net1899),
    .A3(net243),
    .B1(_3649_),
    .X(_1297_));
 sky130_fd_sc_hd__and2_1 _7104_ (.A(net336),
    .B(net244),
    .X(_3650_));
 sky130_fd_sc_hd__a31o_1 _7105_ (.A1(net467),
    .A2(net1806),
    .A3(net242),
    .B1(_3650_),
    .X(_1298_));
 sky130_fd_sc_hd__and2_1 _7106_ (.A(net338),
    .B(net245),
    .X(_3651_));
 sky130_fd_sc_hd__a31o_1 _7107_ (.A1(net443),
    .A2(net1830),
    .A3(net243),
    .B1(_3651_),
    .X(_1299_));
 sky130_fd_sc_hd__and2_1 _7108_ (.A(net337),
    .B(net245),
    .X(_3652_));
 sky130_fd_sc_hd__a31o_1 _7109_ (.A1(net444),
    .A2(net1597),
    .A3(net243),
    .B1(_3652_),
    .X(_1300_));
 sky130_fd_sc_hd__and2_1 _7110_ (.A(net335),
    .B(net244),
    .X(_3653_));
 sky130_fd_sc_hd__a31o_1 _7111_ (.A1(net453),
    .A2(net1858),
    .A3(net242),
    .B1(_3653_),
    .X(_1301_));
 sky130_fd_sc_hd__and2_1 _7112_ (.A(net348),
    .B(net245),
    .X(_3654_));
 sky130_fd_sc_hd__a31o_1 _7113_ (.A1(net440),
    .A2(net1633),
    .A3(net243),
    .B1(_3654_),
    .X(_1302_));
 sky130_fd_sc_hd__and2_1 _7114_ (.A(net346),
    .B(net245),
    .X(_3655_));
 sky130_fd_sc_hd__a31o_1 _7115_ (.A1(net439),
    .A2(net1947),
    .A3(net243),
    .B1(_3655_),
    .X(_1303_));
 sky130_fd_sc_hd__and2_1 _7116_ (.A(net347),
    .B(net245),
    .X(_3656_));
 sky130_fd_sc_hd__a31o_1 _7117_ (.A1(net439),
    .A2(net1409),
    .A3(net243),
    .B1(_3656_),
    .X(_1304_));
 sky130_fd_sc_hd__and2_1 _7118_ (.A(net370),
    .B(net245),
    .X(_3657_));
 sky130_fd_sc_hd__a31o_1 _7119_ (.A1(net446),
    .A2(net1874),
    .A3(net243),
    .B1(_3657_),
    .X(_1305_));
 sky130_fd_sc_hd__nor3_2 _7120_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2758_),
    .Y(_3658_));
 sky130_fd_sc_hd__or3_4 _7121_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2758_),
    .X(_3659_));
 sky130_fd_sc_hd__or3_1 _7122_ (.A(net481),
    .B(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ),
    .C(net240),
    .X(_3660_));
 sky130_fd_sc_hd__o21a_1 _7123_ (.A1(net2046),
    .A2(net238),
    .B1(_3660_),
    .X(_1306_));
 sky130_fd_sc_hd__and2_1 _7124_ (.A(_1679_),
    .B(net240),
    .X(_3661_));
 sky130_fd_sc_hd__a31o_1 _7125_ (.A1(net471),
    .A2(net1750),
    .A3(net238),
    .B1(_3661_),
    .X(_1307_));
 sky130_fd_sc_hd__and2_1 _7126_ (.A(_1667_),
    .B(net240),
    .X(_3662_));
 sky130_fd_sc_hd__a31o_1 _7127_ (.A1(net470),
    .A2(net1792),
    .A3(_3659_),
    .B1(_3662_),
    .X(_1308_));
 sky130_fd_sc_hd__and2_1 _7128_ (.A(_1655_),
    .B(net240),
    .X(_3663_));
 sky130_fd_sc_hd__a31o_1 _7129_ (.A1(net469),
    .A2(net1734),
    .A3(net238),
    .B1(_3663_),
    .X(_1309_));
 sky130_fd_sc_hd__and2_1 _7130_ (.A(_1716_),
    .B(net240),
    .X(_3664_));
 sky130_fd_sc_hd__a31o_1 _7131_ (.A1(net463),
    .A2(net1784),
    .A3(net239),
    .B1(_3664_),
    .X(_1310_));
 sky130_fd_sc_hd__or3b_1 _7132_ (.A(net480),
    .B(net241),
    .C_N(net2146),
    .X(_3665_));
 sky130_fd_sc_hd__o21ai_1 _7133_ (.A1(_1740_),
    .A2(_3659_),
    .B1(_3665_),
    .Y(_1311_));
 sky130_fd_sc_hd__and2_1 _7134_ (.A(_1728_),
    .B(net240),
    .X(_3666_));
 sky130_fd_sc_hd__a31o_1 _7135_ (.A1(net460),
    .A2(net1834),
    .A3(net238),
    .B1(_3666_),
    .X(_1312_));
 sky130_fd_sc_hd__and2_1 _7136_ (.A(net330),
    .B(net241),
    .X(_3667_));
 sky130_fd_sc_hd__a31o_1 _7137_ (.A1(net439),
    .A2(net1746),
    .A3(net239),
    .B1(_3667_),
    .X(_1313_));
 sky130_fd_sc_hd__and2_1 _7138_ (.A(net325),
    .B(net241),
    .X(_3668_));
 sky130_fd_sc_hd__a31o_1 _7139_ (.A1(net448),
    .A2(net1945),
    .A3(net239),
    .B1(_3668_),
    .X(_1314_));
 sky130_fd_sc_hd__and2_1 _7140_ (.A(_1757_),
    .B(net240),
    .X(_3669_));
 sky130_fd_sc_hd__a31o_1 _7141_ (.A1(net460),
    .A2(net1689),
    .A3(net238),
    .B1(_3669_),
    .X(_1315_));
 sky130_fd_sc_hd__and2_1 _7142_ (.A(net326),
    .B(net241),
    .X(_3670_));
 sky130_fd_sc_hd__a31o_1 _7143_ (.A1(net454),
    .A2(net1766),
    .A3(net239),
    .B1(_3670_),
    .X(_1316_));
 sky130_fd_sc_hd__and2_1 _7144_ (.A(net324),
    .B(net241),
    .X(_3671_));
 sky130_fd_sc_hd__a31o_1 _7145_ (.A1(net442),
    .A2(net1629),
    .A3(net239),
    .B1(_3671_),
    .X(_1317_));
 sky130_fd_sc_hd__and2_1 _7146_ (.A(net321),
    .B(net240),
    .X(_3672_));
 sky130_fd_sc_hd__a31o_1 _7147_ (.A1(net463),
    .A2(net1782),
    .A3(net238),
    .B1(_3672_),
    .X(_1318_));
 sky130_fd_sc_hd__and2_1 _7148_ (.A(net323),
    .B(net240),
    .X(_3673_));
 sky130_fd_sc_hd__a31o_1 _7149_ (.A1(net462),
    .A2(net1917),
    .A3(net238),
    .B1(_3673_),
    .X(_1319_));
 sky130_fd_sc_hd__and2_1 _7150_ (.A(_1810_),
    .B(net240),
    .X(_3674_));
 sky130_fd_sc_hd__a31o_1 _7151_ (.A1(net471),
    .A2(net1860),
    .A3(net238),
    .B1(_3674_),
    .X(_1320_));
 sky130_fd_sc_hd__and2_1 _7152_ (.A(net320),
    .B(net240),
    .X(_3675_));
 sky130_fd_sc_hd__a31o_1 _7153_ (.A1(net458),
    .A2(net1846),
    .A3(net238),
    .B1(_3675_),
    .X(_1321_));
 sky130_fd_sc_hd__and2_1 _7154_ (.A(net344),
    .B(net241),
    .X(_3676_));
 sky130_fd_sc_hd__a31o_1 _7155_ (.A1(net452),
    .A2(net1854),
    .A3(net239),
    .B1(_3676_),
    .X(_1322_));
 sky130_fd_sc_hd__nor2_1 _7156_ (.A(_1511_),
    .B(net238),
    .Y(_3677_));
 sky130_fd_sc_hd__a31o_1 _7157_ (.A1(net452),
    .A2(net1893),
    .A3(net238),
    .B1(_3677_),
    .X(_1323_));
 sky130_fd_sc_hd__and2_1 _7158_ (.A(net343),
    .B(net240),
    .X(_3678_));
 sky130_fd_sc_hd__a31o_1 _7159_ (.A1(net465),
    .A2(net1778),
    .A3(net238),
    .B1(_3678_),
    .X(_1324_));
 sky130_fd_sc_hd__and2_1 _7160_ (.A(net345),
    .B(net240),
    .X(_3679_));
 sky130_fd_sc_hd__a31o_1 _7161_ (.A1(net467),
    .A2(net1752),
    .A3(net238),
    .B1(_3679_),
    .X(_1325_));
 sky130_fd_sc_hd__and2_1 _7162_ (.A(net340),
    .B(net241),
    .X(_3680_));
 sky130_fd_sc_hd__a31o_1 _7163_ (.A1(net443),
    .A2(net1762),
    .A3(net239),
    .B1(_3680_),
    .X(_1326_));
 sky130_fd_sc_hd__and2_1 _7164_ (.A(net342),
    .B(net241),
    .X(_3681_));
 sky130_fd_sc_hd__a31o_1 _7165_ (.A1(net444),
    .A2(net1643),
    .A3(net239),
    .B1(_3681_),
    .X(_1327_));
 sky130_fd_sc_hd__and2_1 _7166_ (.A(_1572_),
    .B(net240),
    .X(_3682_));
 sky130_fd_sc_hd__a31o_1 _7167_ (.A1(net467),
    .A2(net1864),
    .A3(net238),
    .B1(_3682_),
    .X(_1328_));
 sky130_fd_sc_hd__and2_1 _7168_ (.A(net339),
    .B(net241),
    .X(_3683_));
 sky130_fd_sc_hd__a31o_1 _7169_ (.A1(net443),
    .A2(net1915),
    .A3(net239),
    .B1(_3683_),
    .X(_1329_));
 sky130_fd_sc_hd__and2_1 _7170_ (.A(_1630_),
    .B(net240),
    .X(_3684_));
 sky130_fd_sc_hd__a31o_1 _7171_ (.A1(net467),
    .A2(net1816),
    .A3(net238),
    .B1(_3684_),
    .X(_1330_));
 sky130_fd_sc_hd__and2_1 _7172_ (.A(net338),
    .B(net241),
    .X(_3685_));
 sky130_fd_sc_hd__a31o_1 _7173_ (.A1(net443),
    .A2(net1836),
    .A3(net239),
    .B1(_3685_),
    .X(_1331_));
 sky130_fd_sc_hd__and2_1 _7174_ (.A(net337),
    .B(net241),
    .X(_3686_));
 sky130_fd_sc_hd__a31o_1 _7175_ (.A1(net444),
    .A2(net1748),
    .A3(net239),
    .B1(_3686_),
    .X(_1332_));
 sky130_fd_sc_hd__and2_1 _7176_ (.A(_1643_),
    .B(net240),
    .X(_3687_));
 sky130_fd_sc_hd__a31o_1 _7177_ (.A1(net453),
    .A2(net1984),
    .A3(net238),
    .B1(_3687_),
    .X(_1333_));
 sky130_fd_sc_hd__and2_1 _7178_ (.A(net348),
    .B(net241),
    .X(_3688_));
 sky130_fd_sc_hd__a31o_1 _7179_ (.A1(net439),
    .A2(net1707),
    .A3(net239),
    .B1(_3688_),
    .X(_1334_));
 sky130_fd_sc_hd__and2_1 _7180_ (.A(net346),
    .B(net241),
    .X(_3689_));
 sky130_fd_sc_hd__a31o_1 _7181_ (.A1(net439),
    .A2(net1722),
    .A3(net239),
    .B1(_3689_),
    .X(_1335_));
 sky130_fd_sc_hd__and2_1 _7182_ (.A(net347),
    .B(net241),
    .X(_3690_));
 sky130_fd_sc_hd__a31o_1 _7183_ (.A1(net439),
    .A2(net1921),
    .A3(net239),
    .B1(_3690_),
    .X(_1336_));
 sky130_fd_sc_hd__and2_1 _7184_ (.A(net370),
    .B(net241),
    .X(_3691_));
 sky130_fd_sc_hd__a31o_1 _7185_ (.A1(net445),
    .A2(net1796),
    .A3(net239),
    .B1(_3691_),
    .X(_1337_));
 sky130_fd_sc_hd__nor2_1 _7186_ (.A(_2266_),
    .B(net163),
    .Y(_1338_));
 sky130_fd_sc_hd__or4_1 _7187_ (.A(net2055),
    .B(net2092),
    .C(net2010),
    .D(_2794_),
    .X(_3692_));
 sky130_fd_sc_hd__a21o_1 _7188_ (.A1(_0066_),
    .A2(_2793_),
    .B1(_2806_),
    .X(_3693_));
 sky130_fd_sc_hd__a2bb2o_1 _7189_ (.A1_N(net2190),
    .A2_N(_2802_),
    .B1(_2803_),
    .B2(_3693_),
    .X(_3694_));
 sky130_fd_sc_hd__a21boi_1 _7190_ (.A1(_2805_),
    .A2(_3694_),
    .B1_N(_2788_),
    .Y(_3695_));
 sky130_fd_sc_hd__o21ai_1 _7191_ (.A1(_2795_),
    .A2(_3695_),
    .B1(net2207),
    .Y(_3696_));
 sky130_fd_sc_hd__o211a_1 _7192_ (.A1(net2190),
    .A2(net2207),
    .B1(_3696_),
    .C1(_2776_),
    .X(_1339_));
 sky130_fd_sc_hd__a211o_1 _7193_ (.A1(net2190),
    .A2(net2010),
    .B1(_2799_),
    .C1(net2092),
    .X(_3697_));
 sky130_fd_sc_hd__a211o_1 _7194_ (.A1(_0067_),
    .A2(_2793_),
    .B1(_2801_),
    .C1(_2806_),
    .X(_3698_));
 sky130_fd_sc_hd__a21bo_1 _7195_ (.A1(_2800_),
    .A2(_3698_),
    .B1_N(_2802_),
    .X(_3699_));
 sky130_fd_sc_hd__a21bo_1 _7196_ (.A1(_3697_),
    .A2(_3699_),
    .B1_N(_2804_),
    .X(_3700_));
 sky130_fd_sc_hd__and3_1 _7197_ (.A(_2776_),
    .B(_2797_),
    .C(_3700_),
    .X(_1340_));
 sky130_fd_sc_hd__a22o_1 _7198_ (.A1(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ),
    .A2(_2801_),
    .B1(_2806_),
    .B2(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .X(_3701_));
 sky130_fd_sc_hd__a31o_1 _7199_ (.A1(_0064_),
    .A2(_2793_),
    .A3(_2807_),
    .B1(_3701_),
    .X(_3702_));
 sky130_fd_sc_hd__nand2_1 _7200_ (.A(_2784_),
    .B(_2790_),
    .Y(_3703_));
 sky130_fd_sc_hd__a32o_1 _7201_ (.A1(_2800_),
    .A2(_3702_),
    .A3(_3703_),
    .B1(_2798_),
    .B2(_2787_),
    .X(_3704_));
 sky130_fd_sc_hd__o211a_1 _7202_ (.A1(net2190),
    .A2(_2802_),
    .B1(_2805_),
    .C1(_3704_),
    .X(_3705_));
 sky130_fd_sc_hd__nor2_1 _7203_ (.A(_2796_),
    .B(_3705_),
    .Y(_3706_));
 sky130_fd_sc_hd__mux2_1 _7204_ (.A0(net2190),
    .A1(_3706_),
    .S(net2207),
    .X(_3707_));
 sky130_fd_sc_hd__nor2_1 _7205_ (.A(net162),
    .B(_3707_),
    .Y(_1341_));
 sky130_fd_sc_hd__nand2_1 _7206_ (.A(net2010),
    .B(_2786_),
    .Y(_3708_));
 sky130_fd_sc_hd__a221o_1 _7207_ (.A1(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .A2(_2785_),
    .B1(_2806_),
    .B2(net2206),
    .C1(_2801_),
    .X(_3709_));
 sky130_fd_sc_hd__a31o_1 _7208_ (.A1(_0065_),
    .A2(_2793_),
    .A3(_2807_),
    .B1(_3709_),
    .X(_3710_));
 sky130_fd_sc_hd__a21bo_1 _7209_ (.A1(_2799_),
    .A2(_3710_),
    .B1_N(_3697_),
    .X(_3711_));
 sky130_fd_sc_hd__a21oi_1 _7210_ (.A1(_3708_),
    .A2(_3711_),
    .B1(_2795_),
    .Y(_3712_));
 sky130_fd_sc_hd__mux2_1 _7211_ (.A0(net2190),
    .A1(_3712_),
    .S(net2207),
    .X(_3713_));
 sky130_fd_sc_hd__nor2_1 _7212_ (.A(net162),
    .B(_3713_),
    .Y(_1342_));
 sky130_fd_sc_hd__and2_1 _7213_ (.A(net468),
    .B(net920),
    .X(_1343_));
 sky130_fd_sc_hd__and2_1 _7214_ (.A(net471),
    .B(net1218),
    .X(_1344_));
 sky130_fd_sc_hd__and2_1 _7215_ (.A(net470),
    .B(net1495),
    .X(_1345_));
 sky130_fd_sc_hd__and2_1 _7216_ (.A(net469),
    .B(net1716),
    .X(_1346_));
 sky130_fd_sc_hd__and2_1 _7217_ (.A(net463),
    .B(net1377),
    .X(_1347_));
 sky130_fd_sc_hd__and2_1 _7218_ (.A(net464),
    .B(net1621),
    .X(_1348_));
 sky130_fd_sc_hd__and2_1 _7219_ (.A(net460),
    .B(net1072),
    .X(_1349_));
 sky130_fd_sc_hd__and2_1 _7220_ (.A(net444),
    .B(net1665),
    .X(_1350_));
 sky130_fd_sc_hd__and2_1 _7221_ (.A(net448),
    .B(net1627),
    .X(_1351_));
 sky130_fd_sc_hd__and2_1 _7222_ (.A(net460),
    .B(net1204),
    .X(_1352_));
 sky130_fd_sc_hd__and2_1 _7223_ (.A(net454),
    .B(net1545),
    .X(_1353_));
 sky130_fd_sc_hd__and2_1 _7224_ (.A(net442),
    .B(net1120),
    .X(_1354_));
 sky130_fd_sc_hd__and2_1 _7225_ (.A(net463),
    .B(net1533),
    .X(_1355_));
 sky130_fd_sc_hd__and2_1 _7226_ (.A(net462),
    .B(net1405),
    .X(_1356_));
 sky130_fd_sc_hd__and2_1 _7227_ (.A(net471),
    .B(net1651),
    .X(_1357_));
 sky130_fd_sc_hd__and2_1 _7228_ (.A(net458),
    .B(net1130),
    .X(_1358_));
 sky130_fd_sc_hd__and2_1 _7229_ (.A(net452),
    .B(net1631),
    .X(_1359_));
 sky130_fd_sc_hd__and2_1 _7230_ (.A(net452),
    .B(net1461),
    .X(_1360_));
 sky130_fd_sc_hd__and2_1 _7231_ (.A(net466),
    .B(net1080),
    .X(_1361_));
 sky130_fd_sc_hd__and2_1 _7232_ (.A(net467),
    .B(net1160),
    .X(_1362_));
 sky130_fd_sc_hd__and2_1 _7233_ (.A(net443),
    .B(net1529),
    .X(_1363_));
 sky130_fd_sc_hd__and2_1 _7234_ (.A(net444),
    .B(net1134),
    .X(_1364_));
 sky130_fd_sc_hd__and2_1 _7235_ (.A(net467),
    .B(net1531),
    .X(_1365_));
 sky130_fd_sc_hd__and2_1 _7236_ (.A(net443),
    .B(net1549),
    .X(_1366_));
 sky130_fd_sc_hd__and2_1 _7237_ (.A(net468),
    .B(net1577),
    .X(_1367_));
 sky130_fd_sc_hd__and2_1 _7238_ (.A(net443),
    .B(net1635),
    .X(_1368_));
 sky130_fd_sc_hd__and2_1 _7239_ (.A(net444),
    .B(net1256),
    .X(_1369_));
 sky130_fd_sc_hd__and2_1 _7240_ (.A(net453),
    .B(net1607),
    .X(_1370_));
 sky130_fd_sc_hd__and2_1 _7241_ (.A(net439),
    .B(net1487),
    .X(_1371_));
 sky130_fd_sc_hd__and2_1 _7242_ (.A(net439),
    .B(net1399),
    .X(_1372_));
 sky130_fd_sc_hd__and2_1 _7243_ (.A(net439),
    .B(net1669),
    .X(_1373_));
 sky130_fd_sc_hd__and2_1 _7244_ (.A(net445),
    .B(net1485),
    .X(_1374_));
 sky130_fd_sc_hd__and3_1 _7245_ (.A(net2019),
    .B(net174),
    .C(net281),
    .X(_1375_));
 sky130_fd_sc_hd__nand2_1 _7246_ (.A(net2019),
    .B(_2265_),
    .Y(_3714_));
 sky130_fd_sc_hd__nand2_1 _7247_ (.A(net2190),
    .B(net2074),
    .Y(_3715_));
 sky130_fd_sc_hd__a21oi_1 _7248_ (.A1(net2020),
    .A2(_3715_),
    .B1(net162),
    .Y(_1376_));
 sky130_fd_sc_hd__nand2_1 _7249_ (.A(net2138),
    .B(net2074),
    .Y(_3716_));
 sky130_fd_sc_hd__a21oi_1 _7250_ (.A1(net2020),
    .A2(_3716_),
    .B1(net162),
    .Y(_1377_));
 sky130_fd_sc_hd__nand2_1 _7251_ (.A(net2007),
    .B(net2074),
    .Y(_3717_));
 sky130_fd_sc_hd__a21oi_1 _7252_ (.A1(net2020),
    .A2(_3717_),
    .B1(net162),
    .Y(_1378_));
 sky130_fd_sc_hd__nand2_1 _7253_ (.A(net2214),
    .B(net2074),
    .Y(_3718_));
 sky130_fd_sc_hd__a21oi_1 _7254_ (.A1(net2020),
    .A2(_3718_),
    .B1(net162),
    .Y(_1379_));
 sky130_fd_sc_hd__nand2_1 _7255_ (.A(net1997),
    .B(_2264_),
    .Y(_3719_));
 sky130_fd_sc_hd__a21oi_1 _7256_ (.A1(net2020),
    .A2(_3719_),
    .B1(net162),
    .Y(_1380_));
 sky130_fd_sc_hd__nand2_1 _7257_ (.A(net1292),
    .B(_2264_),
    .Y(_3720_));
 sky130_fd_sc_hd__a21oi_1 _7258_ (.A1(_3714_),
    .A2(net1293),
    .B1(net162),
    .Y(_1381_));
 sky130_fd_sc_hd__nand2_1 _7259_ (.A(net2172),
    .B(net2074),
    .Y(_3721_));
 sky130_fd_sc_hd__a21oi_1 _7260_ (.A1(net2020),
    .A2(_3721_),
    .B1(net162),
    .Y(_1382_));
 sky130_fd_sc_hd__nand2_1 _7261_ (.A(net381),
    .B(net2074),
    .Y(_3722_));
 sky130_fd_sc_hd__a21oi_1 _7262_ (.A1(net2020),
    .A2(_3722_),
    .B1(net162),
    .Y(_1383_));
 sky130_fd_sc_hd__nand2_1 _7263_ (.A(net385),
    .B(net2074),
    .Y(_3723_));
 sky130_fd_sc_hd__a21oi_1 _7264_ (.A1(net2020),
    .A2(_3723_),
    .B1(net162),
    .Y(_1384_));
 sky130_fd_sc_hd__nand2_1 _7265_ (.A(net392),
    .B(net2074),
    .Y(_3724_));
 sky130_fd_sc_hd__a21oi_1 _7266_ (.A1(net2020),
    .A2(_3724_),
    .B1(net162),
    .Y(_1385_));
 sky130_fd_sc_hd__nand2_1 _7267_ (.A(net402),
    .B(net2074),
    .Y(_3725_));
 sky130_fd_sc_hd__a21oi_1 _7268_ (.A1(net2020),
    .A2(_3725_),
    .B1(net162),
    .Y(_1386_));
 sky130_fd_sc_hd__nand2_1 _7269_ (.A(net2105),
    .B(_2810_),
    .Y(_3726_));
 sky130_fd_sc_hd__nand3_4 _7270_ (.A(net2019),
    .B(net2059),
    .C(_2809_),
    .Y(_3727_));
 sky130_fd_sc_hd__a21oi_1 _7271_ (.A1(net2106),
    .A2(_3727_),
    .B1(net163),
    .Y(_1387_));
 sky130_fd_sc_hd__nand2_1 _7272_ (.A(net409),
    .B(_2810_),
    .Y(_3728_));
 sky130_fd_sc_hd__a21oi_1 _7273_ (.A1(_3727_),
    .A2(_3728_),
    .B1(net163),
    .Y(_1388_));
 sky130_fd_sc_hd__nand2_1 _7274_ (.A(net416),
    .B(_2810_),
    .Y(_3729_));
 sky130_fd_sc_hd__a21oi_1 _7275_ (.A1(_3727_),
    .A2(net2182),
    .B1(net163),
    .Y(_1389_));
 sky130_fd_sc_hd__nand2_1 _7276_ (.A(net426),
    .B(_2810_),
    .Y(_3730_));
 sky130_fd_sc_hd__a21oi_1 _7277_ (.A1(_3727_),
    .A2(net2170),
    .B1(net163),
    .Y(_1390_));
 sky130_fd_sc_hd__nand2_1 _7278_ (.A(net432),
    .B(_2810_),
    .Y(_3731_));
 sky130_fd_sc_hd__a21oi_1 _7279_ (.A1(_3727_),
    .A2(net2144),
    .B1(net163),
    .Y(_1391_));
 sky130_fd_sc_hd__nand2_1 _7280_ (.A(net2055),
    .B(_2810_),
    .Y(_3732_));
 sky130_fd_sc_hd__a21oi_1 _7281_ (.A1(_3727_),
    .A2(net2056),
    .B1(net163),
    .Y(_1392_));
 sky130_fd_sc_hd__nand2_1 _7282_ (.A(net2092),
    .B(_2810_),
    .Y(_3733_));
 sky130_fd_sc_hd__a21oi_1 _7283_ (.A1(_3727_),
    .A2(net2093),
    .B1(net163),
    .Y(_1393_));
 sky130_fd_sc_hd__nand2_1 _7284_ (.A(net2010),
    .B(_2810_),
    .Y(_3734_));
 sky130_fd_sc_hd__a21oi_1 _7285_ (.A1(_3727_),
    .A2(net2011),
    .B1(net163),
    .Y(_1394_));
 sky130_fd_sc_hd__nor2_1 _7286_ (.A(_2790_),
    .B(_3727_),
    .Y(_3735_));
 sky130_fd_sc_hd__a32o_1 _7287_ (.A1(net408),
    .A2(net2058),
    .A3(_2262_),
    .B1(_2790_),
    .B2(net2128),
    .X(_3736_));
 sky130_fd_sc_hd__o21a_1 _7288_ (.A1(_3735_),
    .A2(_3736_),
    .B1(_2776_),
    .X(_1395_));
 sky130_fd_sc_hd__and3_1 _7289_ (.A(net2190),
    .B(net2059),
    .C(_2776_),
    .X(_1396_));
 sky130_fd_sc_hd__and3_1 _7290_ (.A(net2138),
    .B(net2059),
    .C(_2776_),
    .X(_1397_));
 sky130_fd_sc_hd__and3_1 _7291_ (.A(net2007),
    .B(_2265_),
    .C(_2776_),
    .X(_1398_));
 sky130_fd_sc_hd__and3_1 _7292_ (.A(net2214),
    .B(net2059),
    .C(_2776_),
    .X(_1399_));
 sky130_fd_sc_hd__and3_1 _7293_ (.A(net1997),
    .B(_2265_),
    .C(_2776_),
    .X(_1400_));
 sky130_fd_sc_hd__and3_1 _7294_ (.A(net1292),
    .B(net2059),
    .C(_2776_),
    .X(_1401_));
 sky130_fd_sc_hd__nor2_1 _7295_ (.A(_2789_),
    .B(_2810_),
    .Y(_3737_));
 sky130_fd_sc_hd__o21ai_4 _7296_ (.A1(_2264_),
    .A2(_2789_),
    .B1(_2809_),
    .Y(_3738_));
 sky130_fd_sc_hd__a22o_1 _7297_ (.A1(net2199),
    .A2(_2789_),
    .B1(_3738_),
    .B2(net2172),
    .X(_3739_));
 sky130_fd_sc_hd__and3_1 _7298_ (.A(net176),
    .B(net278),
    .C(_3739_),
    .X(_1402_));
 sky130_fd_sc_hd__a22o_1 _7299_ (.A1(net2134),
    .A2(_2789_),
    .B1(_3738_),
    .B2(net382),
    .X(_3740_));
 sky130_fd_sc_hd__and3_1 _7300_ (.A(net2044),
    .B(net286),
    .C(_3740_),
    .X(_1403_));
 sky130_fd_sc_hd__a22o_1 _7301_ (.A1(net2103),
    .A2(_2789_),
    .B1(_3738_),
    .B2(net387),
    .X(_3741_));
 sky130_fd_sc_hd__and3_1 _7302_ (.A(net184),
    .B(net286),
    .C(_3741_),
    .X(_1404_));
 sky130_fd_sc_hd__a22o_1 _7303_ (.A1(net2204),
    .A2(_2789_),
    .B1(_3738_),
    .B2(net398),
    .X(_3742_));
 sky130_fd_sc_hd__and3_1 _7304_ (.A(net179),
    .B(net284),
    .C(_3742_),
    .X(_1405_));
 sky130_fd_sc_hd__a32o_1 _7305_ (.A1(net2128),
    .A2(_1407_),
    .A3(_2789_),
    .B1(_3737_),
    .B2(net408),
    .X(_3743_));
 sky130_fd_sc_hd__and3_1 _7306_ (.A(net176),
    .B(net278),
    .C(_3743_),
    .X(_1406_));
 sky130_fd_sc_hd__o31a_1 _7307_ (.A1(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .A2(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .A3(_2267_),
    .B1(_2266_),
    .X(_3745_));
 sky130_fd_sc_hd__o31a_1 _7308_ (.A1(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .A2(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .A3(_2267_),
    .B1(_2266_),
    .X(_3746_));
 sky130_fd_sc_hd__o31a_1 _7309_ (.A1(net2234),
    .A2(net2203),
    .A3(_2267_),
    .B1(_2266_),
    .X(_3747_));
 sky130_fd_sc_hd__o31a_1 _7310_ (.A1(net2194),
    .A2(net2203),
    .A3(_2267_),
    .B1(_2266_),
    .X(_3748_));
 sky130_fd_sc_hd__inv_2 _7311_ (.A(net480),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _7312_ (.A(net480),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _7313_ (.A(net478),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _7314_ (.A(net476),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _7315_ (.A(net476),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _7316_ (.A(net476),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _7317_ (.A(net478),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _7318_ (.A(net477),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _7319_ (.A(net476),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _7320_ (.A(net476),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _7321_ (.A(net478),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _7322_ (.A(net478),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _7323_ (.A(net478),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _7324_ (.A(net478),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _7325_ (.A(net478),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _7326_ (.A(net480),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _7327_ (.A(net478),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _7328_ (.A(net481),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _7329_ (.A(net474),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _7330_ (.A(net477),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _7331_ (.A(net473),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _7332_ (.A(net477),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _7333_ (.A(net473),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _7334_ (.A(net473),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _7335_ (.A(net473),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _7336_ (.A(net475),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _7337_ (.A(net475),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _7338_ (.A(net475),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _7339_ (.A(net477),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _7340__2 (.A(clknet_leaf_31_clk),
    .Y(net490));
 sky130_fd_sc_hd__inv_2 _7341__3 (.A(clknet_leaf_36_clk),
    .Y(net491));
 sky130_fd_sc_hd__inv_2 _7342__4 (.A(clknet_leaf_32_clk),
    .Y(net492));
 sky130_fd_sc_hd__inv_2 _7343__5 (.A(clknet_leaf_27_clk),
    .Y(net493));
 sky130_fd_sc_hd__inv_2 _7344__6 (.A(clknet_leaf_19_clk),
    .Y(net494));
 sky130_fd_sc_hd__inv_2 _7345__7 (.A(clknet_leaf_44_clk),
    .Y(net495));
 sky130_fd_sc_hd__inv_2 _7346__8 (.A(clknet_leaf_68_clk),
    .Y(net496));
 sky130_fd_sc_hd__inv_2 _7347__9 (.A(clknet_leaf_66_clk),
    .Y(net497));
 sky130_fd_sc_hd__inv_2 _7348__10 (.A(clknet_leaf_45_clk),
    .Y(net498));
 sky130_fd_sc_hd__inv_2 _7349__11 (.A(clknet_leaf_6_clk),
    .Y(net499));
 sky130_fd_sc_hd__inv_2 _7350__12 (.A(clknet_leaf_65_clk),
    .Y(net500));
 sky130_fd_sc_hd__inv_2 _7351__13 (.A(clknet_leaf_46_clk),
    .Y(net501));
 sky130_fd_sc_hd__inv_2 _7352__14 (.A(clknet_leaf_41_clk),
    .Y(net502));
 sky130_fd_sc_hd__inv_2 _7353__15 (.A(clknet_leaf_25_clk),
    .Y(net503));
 sky130_fd_sc_hd__inv_2 _7354__16 (.A(clknet_leaf_10_clk),
    .Y(net504));
 sky130_fd_sc_hd__inv_2 _7355__17 (.A(clknet_leaf_50_clk),
    .Y(net505));
 sky130_fd_sc_hd__inv_2 _7356__18 (.A(clknet_leaf_47_clk),
    .Y(net506));
 sky130_fd_sc_hd__inv_2 _7357__19 (.A(clknet_leaf_25_clk),
    .Y(net507));
 sky130_fd_sc_hd__inv_2 _7358__20 (.A(clknet_leaf_33_clk),
    .Y(net508));
 sky130_fd_sc_hd__inv_2 _7359__21 (.A(clknet_leaf_63_clk),
    .Y(net509));
 sky130_fd_sc_hd__inv_2 _7360__22 (.A(clknet_leaf_59_clk),
    .Y(net510));
 sky130_fd_sc_hd__inv_2 _7361__23 (.A(clknet_leaf_40_clk),
    .Y(net511));
 sky130_fd_sc_hd__inv_2 _7362__24 (.A(clknet_leaf_62_clk),
    .Y(net512));
 sky130_fd_sc_hd__inv_2 _7363__25 (.A(clknet_leaf_46_clk),
    .Y(net513));
 sky130_fd_sc_hd__inv_2 _7364__26 (.A(clknet_leaf_62_clk),
    .Y(net514));
 sky130_fd_sc_hd__inv_2 _7365__27 (.A(clknet_leaf_58_clk),
    .Y(net515));
 sky130_fd_sc_hd__inv_2 _7366__28 (.A(clknet_leaf_51_clk),
    .Y(net516));
 sky130_fd_sc_hd__inv_2 _7367__29 (.A(clknet_leaf_71_clk),
    .Y(net517));
 sky130_fd_sc_hd__inv_2 _7368__30 (.A(clknet_leaf_70_clk),
    .Y(net518));
 sky130_fd_sc_hd__inv_2 _7369__31 (.A(clknet_leaf_70_clk),
    .Y(net519));
 sky130_fd_sc_hd__inv_2 _7370__32 (.A(clknet_leaf_53_clk),
    .Y(net520));
 sky130_fd_sc_hd__inv_2 _7371__33 (.A(clknet_leaf_55_clk),
    .Y(net521));
 sky130_fd_sc_hd__inv_2 _7372__34 (.A(clknet_leaf_2_clk),
    .Y(net522));
 sky130_fd_sc_hd__inv_2 _7373__35 (.A(clknet_leaf_2_clk),
    .Y(net523));
 sky130_fd_sc_hd__inv_2 _7374__36 (.A(clknet_leaf_35_clk),
    .Y(net524));
 sky130_fd_sc_hd__inv_2 _7375__37 (.A(clknet_leaf_34_clk),
    .Y(net525));
 sky130_fd_sc_hd__inv_2 _7376__38 (.A(clknet_leaf_17_clk),
    .Y(net526));
 sky130_fd_sc_hd__inv_2 _7377__39 (.A(clknet_leaf_14_clk),
    .Y(net527));
 sky130_fd_sc_hd__inv_2 _7378__40 (.A(clknet_leaf_56_clk),
    .Y(net528));
 sky130_fd_sc_hd__inv_2 _7379__41 (.A(clknet_leaf_74_clk),
    .Y(net529));
 sky130_fd_sc_hd__inv_2 _7380__42 (.A(clknet_leaf_15_clk),
    .Y(net530));
 sky130_fd_sc_hd__inv_2 _7381__43 (.A(clknet_leaf_35_clk),
    .Y(net531));
 sky130_fd_sc_hd__inv_2 _7382__44 (.A(clknet_leaf_74_clk),
    .Y(net532));
 sky130_fd_sc_hd__inv_2 _7383__45 (.A(clknet_leaf_15_clk),
    .Y(net533));
 sky130_fd_sc_hd__inv_2 _7384__46 (.A(clknet_leaf_56_clk),
    .Y(net534));
 sky130_fd_sc_hd__inv_2 _7385__47 (.A(clknet_leaf_14_clk),
    .Y(net535));
 sky130_fd_sc_hd__inv_2 _7386__48 (.A(clknet_leaf_15_clk),
    .Y(net536));
 sky130_fd_sc_hd__inv_2 _7387__49 (.A(clknet_leaf_14_clk),
    .Y(net537));
 sky130_fd_sc_hd__inv_2 _7388__50 (.A(clknet_leaf_14_clk),
    .Y(net538));
 sky130_fd_sc_hd__inv_2 _7389__51 (.A(clknet_leaf_21_clk),
    .Y(net539));
 sky130_fd_sc_hd__inv_2 _7390__52 (.A(clknet_leaf_14_clk),
    .Y(net540));
 sky130_fd_sc_hd__inv_2 _7391__53 (.A(clknet_leaf_74_clk),
    .Y(net541));
 sky130_fd_sc_hd__inv_2 _7392__54 (.A(clknet_leaf_74_clk),
    .Y(net542));
 sky130_fd_sc_hd__inv_2 _7393__55 (.A(clknet_leaf_18_clk),
    .Y(net543));
 sky130_fd_sc_hd__inv_2 _7394__56 (.A(clknet_leaf_60_clk),
    .Y(net544));
 sky130_fd_sc_hd__inv_2 _7395__57 (.A(clknet_leaf_38_clk),
    .Y(net545));
 sky130_fd_sc_hd__inv_2 _7396__58 (.A(clknet_leaf_52_clk),
    .Y(net546));
 sky130_fd_sc_hd__inv_2 _7397__59 (.A(clknet_leaf_74_clk),
    .Y(net547));
 sky130_fd_sc_hd__inv_2 _7398__60 (.A(clknet_leaf_40_clk),
    .Y(net548));
 sky130_fd_sc_hd__inv_2 _7399__61 (.A(clknet_leaf_74_clk),
    .Y(net549));
 sky130_fd_sc_hd__inv_2 _7400__62 (.A(clknet_leaf_70_clk),
    .Y(net550));
 sky130_fd_sc_hd__inv_2 _7401__63 (.A(clknet_leaf_42_clk),
    .Y(net551));
 sky130_fd_sc_hd__inv_2 _7402__64 (.A(clknet_leaf_57_clk),
    .Y(net552));
 sky130_fd_sc_hd__inv_2 _7403__65 (.A(clknet_leaf_3_clk),
    .Y(net553));
 sky130_fd_sc_hd__inv_2 _7404__66 (.A(clknet_leaf_42_clk),
    .Y(net554));
 sky130_fd_sc_hd__inv_2 _7405__67 (.A(clknet_leaf_42_clk),
    .Y(net555));
 sky130_fd_sc_hd__inv_2 _7406__68 (.A(clknet_leaf_31_clk),
    .Y(net556));
 sky130_fd_sc_hd__inv_2 _7407__69 (.A(clknet_leaf_16_clk),
    .Y(net557));
 sky130_fd_sc_hd__inv_2 _7408__70 (.A(clknet_leaf_10_clk),
    .Y(net558));
 sky130_fd_sc_hd__inv_2 _7409__71 (.A(clknet_leaf_27_clk),
    .Y(net559));
 sky130_fd_sc_hd__inv_2 _7410__72 (.A(clknet_leaf_51_clk),
    .Y(net560));
 sky130_fd_sc_hd__inv_2 _7411__73 (.A(clknet_leaf_62_clk),
    .Y(net561));
 sky130_fd_sc_hd__inv_2 _7412__74 (.A(clknet_leaf_5_clk),
    .Y(net562));
 sky130_fd_sc_hd__inv_2 _7413__75 (.A(clknet_leaf_28_clk),
    .Y(net563));
 sky130_fd_sc_hd__inv_2 _7414__76 (.A(clknet_leaf_4_clk),
    .Y(net564));
 sky130_fd_sc_hd__inv_2 _7415__77 (.A(clknet_leaf_5_clk),
    .Y(net565));
 sky130_fd_sc_hd__inv_2 _7416__78 (.A(clknet_leaf_47_clk),
    .Y(net566));
 sky130_fd_sc_hd__inv_2 _7417__79 (.A(clknet_leaf_45_clk),
    .Y(net567));
 sky130_fd_sc_hd__inv_2 _7418__80 (.A(clknet_leaf_27_clk),
    .Y(net568));
 sky130_fd_sc_hd__inv_2 _7419__81 (.A(clknet_leaf_16_clk),
    .Y(net569));
 sky130_fd_sc_hd__inv_2 _7420__82 (.A(clknet_leaf_51_clk),
    .Y(net570));
 sky130_fd_sc_hd__inv_2 _7421__83 (.A(clknet_leaf_48_clk),
    .Y(net571));
 sky130_fd_sc_hd__inv_2 _7422__84 (.A(clknet_leaf_25_clk),
    .Y(net572));
 sky130_fd_sc_hd__inv_2 _7423__85 (.A(clknet_leaf_24_clk),
    .Y(net573));
 sky130_fd_sc_hd__inv_2 _7424__86 (.A(clknet_leaf_63_clk),
    .Y(net574));
 sky130_fd_sc_hd__inv_2 _7425__87 (.A(clknet_leaf_55_clk),
    .Y(net575));
 sky130_fd_sc_hd__inv_2 _7426__88 (.A(clknet_leaf_40_clk),
    .Y(net576));
 sky130_fd_sc_hd__inv_2 _7427__89 (.A(clknet_leaf_62_clk),
    .Y(net577));
 sky130_fd_sc_hd__inv_2 _7428__90 (.A(clknet_leaf_47_clk),
    .Y(net578));
 sky130_fd_sc_hd__inv_2 _7429__91 (.A(clknet_leaf_62_clk),
    .Y(net579));
 sky130_fd_sc_hd__inv_2 _7430__92 (.A(clknet_leaf_55_clk),
    .Y(net580));
 sky130_fd_sc_hd__inv_2 _7431__93 (.A(clknet_leaf_52_clk),
    .Y(net581));
 sky130_fd_sc_hd__inv_2 _7432__94 (.A(clknet_leaf_0_clk),
    .Y(net582));
 sky130_fd_sc_hd__inv_2 _7433__95 (.A(clknet_leaf_67_clk),
    .Y(net583));
 sky130_fd_sc_hd__inv_2 _7434__96 (.A(clknet_leaf_0_clk),
    .Y(net584));
 sky130_fd_sc_hd__inv_2 _7435__97 (.A(clknet_leaf_52_clk),
    .Y(net585));
 sky130_fd_sc_hd__inv_2 _7436__98 (.A(clknet_leaf_36_clk),
    .Y(net586));
 sky130_fd_sc_hd__inv_2 _7437__99 (.A(clknet_leaf_31_clk),
    .Y(net587));
 sky130_fd_sc_hd__inv_2 _7438__100 (.A(clknet_leaf_36_clk),
    .Y(net588));
 sky130_fd_sc_hd__inv_2 _7439__101 (.A(clknet_leaf_24_clk),
    .Y(net589));
 sky130_fd_sc_hd__inv_2 _7440__102 (.A(clknet_leaf_29_clk),
    .Y(net590));
 sky130_fd_sc_hd__inv_2 _7441__103 (.A(clknet_leaf_25_clk),
    .Y(net591));
 sky130_fd_sc_hd__inv_2 _7442__104 (.A(clknet_leaf_44_clk),
    .Y(net592));
 sky130_fd_sc_hd__inv_2 _7443__105 (.A(clknet_leaf_68_clk),
    .Y(net593));
 sky130_fd_sc_hd__inv_2 _7444__106 (.A(clknet_leaf_5_clk),
    .Y(net594));
 sky130_fd_sc_hd__inv_2 _7445__107 (.A(clknet_leaf_44_clk),
    .Y(net595));
 sky130_fd_sc_hd__inv_2 _7446__108 (.A(clknet_leaf_6_clk),
    .Y(net596));
 sky130_fd_sc_hd__inv_2 _7447__109 (.A(clknet_leaf_65_clk),
    .Y(net597));
 sky130_fd_sc_hd__inv_2 _7448__110 (.A(clknet_leaf_30_clk),
    .Y(net598));
 sky130_fd_sc_hd__inv_2 _7449__111 (.A(clknet_leaf_45_clk),
    .Y(net599));
 sky130_fd_sc_hd__inv_2 _7450__112 (.A(clknet_leaf_25_clk),
    .Y(net600));
 sky130_fd_sc_hd__inv_2 _7451__113 (.A(clknet_leaf_10_clk),
    .Y(net601));
 sky130_fd_sc_hd__inv_2 _7452__114 (.A(clknet_leaf_48_clk),
    .Y(net602));
 sky130_fd_sc_hd__inv_2 _7453__115 (.A(clknet_leaf_47_clk),
    .Y(net603));
 sky130_fd_sc_hd__inv_2 _7454__116 (.A(clknet_leaf_25_clk),
    .Y(net604));
 sky130_fd_sc_hd__inv_2 _7455__117 (.A(clknet_leaf_33_clk),
    .Y(net605));
 sky130_fd_sc_hd__inv_2 _7456__118 (.A(clknet_leaf_59_clk),
    .Y(net606));
 sky130_fd_sc_hd__inv_2 _7457__119 (.A(clknet_leaf_58_clk),
    .Y(net607));
 sky130_fd_sc_hd__inv_2 _7458__120 (.A(clknet_leaf_40_clk),
    .Y(net608));
 sky130_fd_sc_hd__inv_2 _7459__121 (.A(clknet_leaf_62_clk),
    .Y(net609));
 sky130_fd_sc_hd__inv_2 _7460__122 (.A(clknet_leaf_46_clk),
    .Y(net610));
 sky130_fd_sc_hd__inv_2 _7461__123 (.A(clknet_leaf_62_clk),
    .Y(net611));
 sky130_fd_sc_hd__inv_2 _7462__124 (.A(clknet_leaf_58_clk),
    .Y(net612));
 sky130_fd_sc_hd__inv_2 _7463__125 (.A(clknet_leaf_51_clk),
    .Y(net613));
 sky130_fd_sc_hd__inv_2 _7464__126 (.A(clknet_leaf_71_clk),
    .Y(net614));
 sky130_fd_sc_hd__inv_2 _7465__127 (.A(clknet_leaf_67_clk),
    .Y(net615));
 sky130_fd_sc_hd__inv_2 _7466__128 (.A(clknet_leaf_66_clk),
    .Y(net616));
 sky130_fd_sc_hd__inv_2 _7467__129 (.A(clknet_leaf_53_clk),
    .Y(net617));
 sky130_fd_sc_hd__inv_2 _7468_ (.A(net480),
    .Y(_0260_));
 sky130_fd_sc_hd__inv_2 _7469_ (.A(net480),
    .Y(_0261_));
 sky130_fd_sc_hd__inv_2 _7470_ (.A(net480),
    .Y(_0262_));
 sky130_fd_sc_hd__inv_2 _7471_ (.A(net478),
    .Y(_0263_));
 sky130_fd_sc_hd__inv_2 _7472_ (.A(net476),
    .Y(_0264_));
 sky130_fd_sc_hd__inv_2 _7473_ (.A(net476),
    .Y(_0265_));
 sky130_fd_sc_hd__inv_2 _7474_ (.A(net476),
    .Y(_0266_));
 sky130_fd_sc_hd__inv_2 _7475_ (.A(net478),
    .Y(_0267_));
 sky130_fd_sc_hd__inv_2 _7476_ (.A(net477),
    .Y(_0268_));
 sky130_fd_sc_hd__inv_2 _7477_ (.A(net476),
    .Y(_0269_));
 sky130_fd_sc_hd__inv_2 _7478_ (.A(net476),
    .Y(_0270_));
 sky130_fd_sc_hd__inv_2 _7479_ (.A(net476),
    .Y(_0271_));
 sky130_fd_sc_hd__inv_2 _7480_ (.A(net478),
    .Y(_0272_));
 sky130_fd_sc_hd__inv_2 _7481_ (.A(net479),
    .Y(_0273_));
 sky130_fd_sc_hd__inv_2 _7482_ (.A(net478),
    .Y(_0274_));
 sky130_fd_sc_hd__inv_2 _7483_ (.A(net479),
    .Y(_0275_));
 sky130_fd_sc_hd__inv_2 _7484_ (.A(net480),
    .Y(_0276_));
 sky130_fd_sc_hd__inv_2 _7485_ (.A(net480),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_2 _7486_ (.A(net480),
    .Y(_0278_));
 sky130_fd_sc_hd__inv_2 _7487_ (.A(net474),
    .Y(_0279_));
 sky130_fd_sc_hd__inv_2 _7488_ (.A(net474),
    .Y(_0280_));
 sky130_fd_sc_hd__inv_2 _7489_ (.A(net474),
    .Y(_0281_));
 sky130_fd_sc_hd__inv_2 _7490_ (.A(net473),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_2 _7491_ (.A(net473),
    .Y(_0283_));
 sky130_fd_sc_hd__inv_2 _7492_ (.A(net473),
    .Y(_0284_));
 sky130_fd_sc_hd__inv_2 _7493_ (.A(net474),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_2 _7494_ (.A(net475),
    .Y(_0286_));
 sky130_fd_sc_hd__inv_2 _7495_ (.A(net475),
    .Y(_0287_));
 sky130_fd_sc_hd__inv_2 _7496_ (.A(net475),
    .Y(_0288_));
 sky130_fd_sc_hd__inv_2 _7497_ (.A(net474),
    .Y(_0289_));
 sky130_fd_sc_hd__dfxtp_4 _7498_ (.CLK(clknet_leaf_51_clk),
    .D(net790),
    .Q(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7499_ (.CLK(clknet_leaf_12_clk),
    .D(net716),
    .Q(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7500_ (.CLK(clknet_leaf_23_clk),
    .D(_0292_),
    .RESET_B(net465),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_4 _7501_ (.CLK(clknet_leaf_19_clk),
    .D(_0293_),
    .RESET_B(_0102_),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_4 _7502_ (.CLK(clknet_leaf_16_clk),
    .D(_0294_),
    .RESET_B(_0103_),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_4 _7503_ (.CLK(clknet_leaf_11_clk),
    .D(_0295_),
    .RESET_B(_0104_),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_4 _7504_ (.CLK(clknet_leaf_9_clk),
    .D(_0296_),
    .RESET_B(_0105_),
    .Q(net126));
 sky130_fd_sc_hd__dfrtp_4 _7505_ (.CLK(clknet_leaf_11_clk),
    .D(_0297_),
    .RESET_B(_0106_),
    .Q(net127));
 sky130_fd_sc_hd__dfrtp_4 _7506_ (.CLK(clknet_leaf_13_clk),
    .D(_0298_),
    .RESET_B(_0107_),
    .Q(net128));
 sky130_fd_sc_hd__dfrtp_4 _7507_ (.CLK(clknet_leaf_9_clk),
    .D(_0299_),
    .RESET_B(_0108_),
    .Q(net129));
 sky130_fd_sc_hd__dfrtp_4 _7508_ (.CLK(clknet_leaf_4_clk),
    .D(_0300_),
    .RESET_B(_0109_),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_4 _7509_ (.CLK(clknet_leaf_13_clk),
    .D(_0301_),
    .RESET_B(_0110_),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_4 _7510_ (.CLK(clknet_leaf_13_clk),
    .D(_0302_),
    .RESET_B(_0111_),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_4 _7511_ (.CLK(clknet_leaf_11_clk),
    .D(_0303_),
    .RESET_B(_0112_),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_4 _7512_ (.CLK(clknet_leaf_15_clk),
    .D(_0304_),
    .RESET_B(_0113_),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_4 _7513_ (.CLK(clknet_leaf_15_clk),
    .D(_0305_),
    .RESET_B(_0114_),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_4 _7514_ (.CLK(clknet_leaf_10_clk),
    .D(_0306_),
    .RESET_B(_0115_),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_4 _7515_ (.CLK(clknet_leaf_10_clk),
    .D(_0307_),
    .RESET_B(_0116_),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_4 _7516_ (.CLK(clknet_leaf_21_clk),
    .D(_0308_),
    .RESET_B(_0117_),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_4 _7517_ (.CLK(clknet_leaf_27_clk),
    .D(_0309_),
    .RESET_B(_0118_),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_4 _7518_ (.CLK(clknet_leaf_32_clk),
    .D(_0310_),
    .RESET_B(_0119_),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_4 _7519_ (.CLK(clknet_leaf_54_clk),
    .D(_0311_),
    .RESET_B(_0120_),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_4 _7520_ (.CLK(clknet_leaf_44_clk),
    .D(_0312_),
    .RESET_B(_0121_),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_4 _7521_ (.CLK(clknet_leaf_58_clk),
    .D(_0313_),
    .RESET_B(_0122_),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_2 _7522_ (.CLK(clknet_leaf_49_clk),
    .D(_0314_),
    .RESET_B(_0123_),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_4 _7523_ (.CLK(clknet_leaf_58_clk),
    .D(_0315_),
    .RESET_B(_0124_),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_2 _7524_ (.CLK(clknet_leaf_58_clk),
    .D(_0316_),
    .RESET_B(_0125_),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_4 _7525_ (.CLK(clknet_leaf_49_clk),
    .D(_0317_),
    .RESET_B(_0126_),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_4 _7526_ (.CLK(clknet_leaf_0_clk),
    .D(_0318_),
    .RESET_B(_0127_),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_4 _7527_ (.CLK(clknet_leaf_74_clk),
    .D(_0319_),
    .RESET_B(_0128_),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_4 _7528_ (.CLK(clknet_leaf_0_clk),
    .D(_0320_),
    .RESET_B(_0129_),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_4 _7529_ (.CLK(clknet_leaf_49_clk),
    .D(_0321_),
    .RESET_B(_0130_),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_1 _7530_ (.CLK(clknet_leaf_23_clk),
    .D(net2132),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7531_ (.CLK(clknet_leaf_16_clk),
    .D(_0323_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7532_ (.CLK(clknet_leaf_19_clk),
    .D(_0324_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7533_ (.CLK(clknet_leaf_13_clk),
    .D(net2006),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7534_ (.CLK(clknet_leaf_9_clk),
    .D(net1983),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7535_ (.CLK(clknet_leaf_9_clk),
    .D(_0327_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7536_ (.CLK(clknet_leaf_13_clk),
    .D(_0328_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7537_ (.CLK(clknet_leaf_9_clk),
    .D(net2002),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7538_ (.CLK(clknet_leaf_3_clk),
    .D(_0330_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7539_ (.CLK(clknet_leaf_3_clk),
    .D(_0331_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7540_ (.CLK(clknet_leaf_3_clk),
    .D(net1950),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7541_ (.CLK(clknet_leaf_11_clk),
    .D(_0333_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7542_ (.CLK(clknet_leaf_15_clk),
    .D(_0334_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7543_ (.CLK(clknet_leaf_15_clk),
    .D(_0335_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7544_ (.CLK(clknet_leaf_10_clk),
    .D(_0336_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7545_ (.CLK(clknet_leaf_10_clk),
    .D(_0337_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7546_ (.CLK(clknet_leaf_21_clk),
    .D(_0338_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7547_ (.CLK(clknet_leaf_27_clk),
    .D(net1334),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7548_ (.CLK(clknet_leaf_34_clk),
    .D(net736),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7549_ (.CLK(clknet_leaf_53_clk),
    .D(net1829),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7550_ (.CLK(clknet_leaf_49_clk),
    .D(_0342_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7551_ (.CLK(clknet_leaf_54_clk),
    .D(net662),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7552_ (.CLK(clknet_leaf_50_clk),
    .D(_0344_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7553_ (.CLK(clknet_leaf_58_clk),
    .D(_0345_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7554_ (.CLK(clknet_leaf_58_clk),
    .D(_0346_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7555_ (.CLK(clknet_leaf_54_clk),
    .D(_0347_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7556_ (.CLK(clknet_leaf_0_clk),
    .D(_0348_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7557_ (.CLK(clknet_leaf_0_clk),
    .D(_0349_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7558_ (.CLK(clknet_leaf_0_clk),
    .D(_0350_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7559_ (.CLK(clknet_leaf_53_clk),
    .D(net1851),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7560_ (.CLK(clknet_leaf_6_clk),
    .D(_0352_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7561_ (.CLK(clknet_leaf_4_clk),
    .D(_0353_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7562_ (.CLK(clknet_leaf_3_clk),
    .D(_0354_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7563_ (.CLK(clknet_leaf_3_clk),
    .D(_0355_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7564_ (.CLK(clknet_leaf_4_clk),
    .D(_0356_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7565_ (.CLK(clknet_leaf_18_clk),
    .D(_0357_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7566_ (.CLK(clknet_leaf_13_clk),
    .D(_0358_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7567_ (.CLK(clknet_leaf_39_clk),
    .D(_0359_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7568_ (.CLK(clknet_leaf_18_clk),
    .D(_0360_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7569_ (.CLK(clknet_leaf_3_clk),
    .D(_0361_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[11] ));
 sky130_fd_sc_hd__dfxtp_2 _7570_ (.CLK(clknet_leaf_52_clk),
    .D(_0362_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7571_ (.CLK(clknet_leaf_18_clk),
    .D(_0363_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7572_ (.CLK(clknet_leaf_21_clk),
    .D(_0364_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__dfxtp_4 _7573_ (.CLK(clknet_leaf_21_clk),
    .D(_0365_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7574_ (.CLK(clknet_leaf_52_clk),
    .D(_0366_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7575_ (.CLK(clknet_leaf_62_clk),
    .D(_0367_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ));
 sky130_fd_sc_hd__dfxtp_4 _7576_ (.CLK(clknet_leaf_71_clk),
    .D(_0368_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7577_ (.CLK(clknet_leaf_39_clk),
    .D(_0369_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[19] ));
 sky130_fd_sc_hd__dfxtp_4 _7578_ (.CLK(clknet_leaf_39_clk),
    .D(_0370_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7579_ (.CLK(clknet_leaf_53_clk),
    .D(_0371_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7580_ (.CLK(clknet_leaf_39_clk),
    .D(_0372_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7581_ (.CLK(clknet_leaf_55_clk),
    .D(_0373_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7582_ (.CLK(clknet_leaf_42_clk),
    .D(_0374_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7583_ (.CLK(clknet_leaf_3_clk),
    .D(_0375_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7584_ (.CLK(clknet_leaf_67_clk),
    .D(_0376_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[26] ));
 sky130_fd_sc_hd__dfxtp_2 _7585_ (.CLK(clknet_leaf_39_clk),
    .D(_0377_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7586_ (.CLK(clknet_leaf_72_clk),
    .D(_0378_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7587_ (.CLK(clknet_leaf_21_clk),
    .D(_0379_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7588_ (.CLK(clknet_leaf_55_clk),
    .D(_0380_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ));
 sky130_fd_sc_hd__dfxtp_1 _7589_ (.CLK(clknet_leaf_3_clk),
    .D(_0381_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7590_ (.CLK(clknet_leaf_24_clk),
    .D(_0382_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7591_ (.CLK(clknet_leaf_25_clk),
    .D(_0383_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7592_ (.CLK(clknet_leaf_28_clk),
    .D(_0384_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7593_ (.CLK(clknet_leaf_11_clk),
    .D(_0385_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7594_ (.CLK(clknet_leaf_8_clk),
    .D(_0386_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7595_ (.CLK(clknet_leaf_12_clk),
    .D(_0387_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7596_ (.CLK(clknet_leaf_1_clk),
    .D(_0388_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7597_ (.CLK(clknet_leaf_8_clk),
    .D(_0389_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7598_ (.CLK(clknet_leaf_4_clk),
    .D(_0390_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7599_ (.CLK(clknet_leaf_12_clk),
    .D(_0391_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7600_ (.CLK(clknet_leaf_15_clk),
    .D(_0392_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7601_ (.CLK(clknet_leaf_9_clk),
    .D(_0393_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7602_ (.CLK(clknet_leaf_10_clk),
    .D(_0394_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7603_ (.CLK(clknet_leaf_16_clk),
    .D(_0395_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7604_ (.CLK(clknet_leaf_11_clk),
    .D(_0396_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7605_ (.CLK(clknet_leaf_27_clk),
    .D(_0397_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7606_ (.CLK(clknet_leaf_21_clk),
    .D(_0398_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7607_ (.CLK(clknet_leaf_27_clk),
    .D(_0399_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7608_ (.CLK(clknet_leaf_58_clk),
    .D(_0400_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7609_ (.CLK(clknet_leaf_53_clk),
    .D(_0401_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7610_ (.CLK(clknet_leaf_44_clk),
    .D(_0402_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7611_ (.CLK(clknet_leaf_63_clk),
    .D(_0403_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7612_ (.CLK(clknet_leaf_50_clk),
    .D(_0404_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7613_ (.CLK(clknet_leaf_58_clk),
    .D(_0405_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7614_ (.CLK(clknet_leaf_58_clk),
    .D(_0406_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7615_ (.CLK(clknet_leaf_48_clk),
    .D(_0407_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7616_ (.CLK(clknet_leaf_66_clk),
    .D(_0408_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7617_ (.CLK(clknet_leaf_0_clk),
    .D(_0409_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7618_ (.CLK(clknet_leaf_65_clk),
    .D(_0410_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7619_ (.CLK(clknet_leaf_49_clk),
    .D(_0411_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7620_ (.CLK(clknet_leaf_35_clk),
    .D(net1696),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7621_ (.CLK(clknet_leaf_35_clk),
    .D(net1195),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7622_ (.CLK(clknet_leaf_35_clk),
    .D(net901),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7623_ (.CLK(clknet_leaf_35_clk),
    .D(net893),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7624_ (.CLK(clknet_leaf_29_clk),
    .D(net1155),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7625_ (.CLK(clknet_leaf_20_clk),
    .D(net1149),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7626_ (.CLK(clknet_leaf_44_clk),
    .D(net1725),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7627_ (.CLK(clknet_leaf_68_clk),
    .D(net1063),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7628_ (.CLK(clknet_leaf_66_clk),
    .D(net1271),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7629_ (.CLK(clknet_leaf_45_clk),
    .D(net1031),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7630_ (.CLK(clknet_leaf_65_clk),
    .D(net1560),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7631_ (.CLK(clknet_leaf_71_clk),
    .D(net1624),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7632_ (.CLK(clknet_leaf_30_clk),
    .D(net1143),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7633_ (.CLK(clknet_leaf_41_clk),
    .D(net1574),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7634_ (.CLK(clknet_leaf_23_clk),
    .D(net1458),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7635_ (.CLK(clknet_leaf_25_clk),
    .D(net1600),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7636_ (.CLK(clknet_leaf_50_clk),
    .D(net1071),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7637_ (.CLK(clknet_leaf_44_clk),
    .D(net1713),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7638_ (.CLK(clknet_leaf_22_clk),
    .D(net1504),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7639_ (.CLK(clknet_leaf_33_clk),
    .D(net1033),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7640_ (.CLK(clknet_leaf_59_clk),
    .D(net1085),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7641_ (.CLK(clknet_leaf_57_clk),
    .D(net969),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7642_ (.CLK(clknet_leaf_40_clk),
    .D(net1694),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7643_ (.CLK(clknet_leaf_62_clk),
    .D(net1642),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7644_ (.CLK(clknet_leaf_40_clk),
    .D(net1510),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7645_ (.CLK(clknet_leaf_61_clk),
    .D(net1604),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7646_ (.CLK(clknet_leaf_57_clk),
    .D(net1187),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7647_ (.CLK(clknet_leaf_50_clk),
    .D(net1528),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7648_ (.CLK(clknet_leaf_70_clk),
    .D(net1626),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7649_ (.CLK(clknet_leaf_69_clk),
    .D(net1103),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7650_ (.CLK(clknet_leaf_70_clk),
    .D(net1326),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7651_ (.CLK(clknet_leaf_54_clk),
    .D(net1041),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7652_ (.CLK(clknet_leaf_36_clk),
    .D(net991),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7653_ (.CLK(clknet_leaf_36_clk),
    .D(net909),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7654_ (.CLK(clknet_leaf_36_clk),
    .D(net1674),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7655_ (.CLK(clknet_leaf_33_clk),
    .D(net1139),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7656_ (.CLK(clknet_leaf_29_clk),
    .D(net1247),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7657_ (.CLK(clknet_leaf_19_clk),
    .D(net1151),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7658_ (.CLK(clknet_leaf_44_clk),
    .D(net1612),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7659_ (.CLK(clknet_leaf_67_clk),
    .D(net1452),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7660_ (.CLK(clknet_leaf_66_clk),
    .D(net1075),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7661_ (.CLK(clknet_leaf_45_clk),
    .D(net1253),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7662_ (.CLK(clknet_leaf_5_clk),
    .D(net1245),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7663_ (.CLK(clknet_leaf_71_clk),
    .D(net1263),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7664_ (.CLK(clknet_leaf_29_clk),
    .D(net1402),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7665_ (.CLK(clknet_leaf_45_clk),
    .D(net1217),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7666_ (.CLK(clknet_leaf_25_clk),
    .D(net1542),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7667_ (.CLK(clknet_leaf_26_clk),
    .D(net1169),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7668_ (.CLK(clknet_leaf_50_clk),
    .D(net1221),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7669_ (.CLK(clknet_leaf_47_clk),
    .D(net1354),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7670_ (.CLK(clknet_leaf_19_clk),
    .D(net1105),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7671_ (.CLK(clknet_leaf_24_clk),
    .D(net1111),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7672_ (.CLK(clknet_leaf_60_clk),
    .D(net997),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7673_ (.CLK(clknet_leaf_57_clk),
    .D(net1025),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7674_ (.CLK(clknet_leaf_37_clk),
    .D(net1185),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7675_ (.CLK(clknet_leaf_62_clk),
    .D(net1552),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7676_ (.CLK(clknet_leaf_46_clk),
    .D(net1047),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7677_ (.CLK(clknet_leaf_69_clk),
    .D(net1302),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7678_ (.CLK(clknet_leaf_60_clk),
    .D(net985),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7679_ (.CLK(clknet_leaf_50_clk),
    .D(net1259),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7680_ (.CLK(clknet_leaf_70_clk),
    .D(net1404),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7681_ (.CLK(clknet_leaf_69_clk),
    .D(net1043),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7682_ (.CLK(clknet_leaf_70_clk),
    .D(net1432),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7683_ (.CLK(clknet_leaf_58_clk),
    .D(net1646),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7684_ (.CLK(clknet_leaf_36_clk),
    .D(net856),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7685_ (.CLK(clknet_leaf_36_clk),
    .D(net1281),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7686_ (.CLK(clknet_leaf_37_clk),
    .D(net1394),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7687_ (.CLK(clknet_leaf_31_clk),
    .D(net862),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7688_ (.CLK(clknet_leaf_29_clk),
    .D(net1330),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7689_ (.CLK(clknet_leaf_25_clk),
    .D(net1566),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7690_ (.CLK(clknet_leaf_44_clk),
    .D(net1698),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7691_ (.CLK(clknet_leaf_68_clk),
    .D(net1091),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7692_ (.CLK(clknet_leaf_67_clk),
    .D(net949),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7693_ (.CLK(clknet_leaf_41_clk),
    .D(net1514),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7694_ (.CLK(clknet_leaf_65_clk),
    .D(net1602),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7695_ (.CLK(clknet_leaf_67_clk),
    .D(net935),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7696_ (.CLK(clknet_leaf_30_clk),
    .D(net1737),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7697_ (.CLK(clknet_leaf_41_clk),
    .D(net1314),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7698_ (.CLK(clknet_leaf_24_clk),
    .D(net1576),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7699_ (.CLK(clknet_leaf_26_clk),
    .D(net1125),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7700_ (.CLK(clknet_leaf_50_clk),
    .D(net1502),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7701_ (.CLK(clknet_leaf_44_clk),
    .D(net1757),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7702_ (.CLK(clknet_leaf_25_clk),
    .D(net1664),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7703_ (.CLK(clknet_leaf_32_clk),
    .D(net1203),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7704_ (.CLK(clknet_leaf_59_clk),
    .D(net1249),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7705_ (.CLK(clknet_leaf_57_clk),
    .D(net1177),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7706_ (.CLK(clknet_leaf_40_clk),
    .D(net1442),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7707_ (.CLK(clknet_leaf_61_clk),
    .D(net1189),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7708_ (.CLK(clknet_leaf_41_clk),
    .D(net1727),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7709_ (.CLK(clknet_leaf_61_clk),
    .D(net1416),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7710_ (.CLK(clknet_leaf_59_clk),
    .D(net1079),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7711_ (.CLK(clknet_leaf_50_clk),
    .D(net1289),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7712_ (.CLK(clknet_leaf_70_clk),
    .D(net1261),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7713_ (.CLK(clknet_leaf_61_clk),
    .D(net1362),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7714_ (.CLK(clknet_leaf_70_clk),
    .D(net1620),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7715_ (.CLK(clknet_leaf_54_clk),
    .D(net1306),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7716_ (.CLK(net489),
    .D(_0000_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7717_ (.CLK(net490),
    .D(_0011_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7718_ (.CLK(net491),
    .D(_0022_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7719_ (.CLK(net492),
    .D(_0025_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7720_ (.CLK(net493),
    .D(_0026_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7721_ (.CLK(net494),
    .D(_0027_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7722_ (.CLK(net495),
    .D(_0028_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7723_ (.CLK(net496),
    .D(_0029_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7724_ (.CLK(net497),
    .D(_0030_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7725_ (.CLK(net498),
    .D(_0031_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7726_ (.CLK(net499),
    .D(_0001_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7727_ (.CLK(net500),
    .D(_0002_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7728_ (.CLK(net501),
    .D(_0003_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7729_ (.CLK(net502),
    .D(_0004_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7730_ (.CLK(net503),
    .D(_0005_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7731_ (.CLK(net504),
    .D(_0006_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7732_ (.CLK(net505),
    .D(_0007_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7733_ (.CLK(net506),
    .D(_0008_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7734_ (.CLK(net507),
    .D(_0009_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7735_ (.CLK(net508),
    .D(_0010_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7736_ (.CLK(net509),
    .D(_0012_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7737_ (.CLK(net510),
    .D(_0013_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7738_ (.CLK(net511),
    .D(_0014_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7739_ (.CLK(net512),
    .D(_0015_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7740_ (.CLK(net513),
    .D(_0016_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7741_ (.CLK(net514),
    .D(_0017_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7742_ (.CLK(net515),
    .D(_0018_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7743_ (.CLK(net516),
    .D(_0019_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7744_ (.CLK(net517),
    .D(_0020_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7745_ (.CLK(net518),
    .D(_0021_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7746_ (.CLK(net519),
    .D(_0023_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7747_ (.CLK(net520),
    .D(_0024_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7748_ (.CLK(clknet_leaf_36_clk),
    .D(net1265),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7749_ (.CLK(clknet_leaf_34_clk),
    .D(net905),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7750_ (.CLK(clknet_leaf_34_clk),
    .D(net983),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7751_ (.CLK(clknet_leaf_35_clk),
    .D(net971),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7752_ (.CLK(clknet_leaf_29_clk),
    .D(net1434),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7753_ (.CLK(clknet_leaf_20_clk),
    .D(net1237),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7754_ (.CLK(clknet_leaf_44_clk),
    .D(net1654),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7755_ (.CLK(clknet_leaf_67_clk),
    .D(net1564),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7756_ (.CLK(clknet_leaf_71_clk),
    .D(net1498),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7757_ (.CLK(clknet_leaf_45_clk),
    .D(net1145),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7758_ (.CLK(clknet_leaf_5_clk),
    .D(net1255),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7759_ (.CLK(clknet_leaf_71_clk),
    .D(net1562),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7760_ (.CLK(clknet_leaf_30_clk),
    .D(net941),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7761_ (.CLK(clknet_leaf_41_clk),
    .D(net1592),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7762_ (.CLK(clknet_leaf_23_clk),
    .D(net1350),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7763_ (.CLK(clknet_leaf_26_clk),
    .D(net1191),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7764_ (.CLK(clknet_leaf_50_clk),
    .D(net1448),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7765_ (.CLK(clknet_leaf_47_clk),
    .D(net1556),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7766_ (.CLK(clknet_leaf_20_clk),
    .D(net1037),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7767_ (.CLK(clknet_leaf_24_clk),
    .D(net1478),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7768_ (.CLK(clknet_leaf_59_clk),
    .D(net1304),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7769_ (.CLK(clknet_leaf_57_clk),
    .D(net1009),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7770_ (.CLK(clknet_leaf_37_clk),
    .D(net1199),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7771_ (.CLK(clknet_leaf_62_clk),
    .D(net1538),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7772_ (.CLK(clknet_leaf_37_clk),
    .D(net1398),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7773_ (.CLK(clknet_leaf_69_clk),
    .D(net1065),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7774_ (.CLK(clknet_leaf_59_clk),
    .D(net1083),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7775_ (.CLK(clknet_leaf_50_clk),
    .D(net1580),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7776_ (.CLK(clknet_leaf_71_clk),
    .D(net1251),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7777_ (.CLK(clknet_leaf_68_clk),
    .D(net1440),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7778_ (.CLK(clknet_leaf_71_clk),
    .D(net1616),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7779_ (.CLK(clknet_leaf_54_clk),
    .D(net1239),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7780_ (.CLK(clknet_leaf_35_clk),
    .D(net1843),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7781_ (.CLK(clknet_leaf_34_clk),
    .D(net867),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7782_ (.CLK(clknet_leaf_35_clk),
    .D(net915),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7783_ (.CLK(clknet_leaf_35_clk),
    .D(net873),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7784_ (.CLK(clknet_leaf_29_clk),
    .D(net1229),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7785_ (.CLK(clknet_leaf_20_clk),
    .D(net931),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7786_ (.CLK(clknet_leaf_44_clk),
    .D(net1360),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7787_ (.CLK(clknet_leaf_67_clk),
    .D(net1061),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7788_ (.CLK(clknet_leaf_71_clk),
    .D(net1207),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7789_ (.CLK(clknet_leaf_45_clk),
    .D(net1167),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7790_ (.CLK(clknet_leaf_5_clk),
    .D(net1183),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7791_ (.CLK(clknet_leaf_71_clk),
    .D(net1456),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7792_ (.CLK(clknet_leaf_30_clk),
    .D(net1001),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7793_ (.CLK(clknet_leaf_41_clk),
    .D(net1490),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7794_ (.CLK(clknet_leaf_23_clk),
    .D(net1243),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7795_ (.CLK(clknet_leaf_25_clk),
    .D(net1805),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7796_ (.CLK(clknet_leaf_50_clk),
    .D(net1733),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7797_ (.CLK(clknet_leaf_47_clk),
    .D(net1175),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7798_ (.CLK(clknet_leaf_21_clk),
    .D(net1338),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7799_ (.CLK(clknet_leaf_24_clk),
    .D(net1320),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7800_ (.CLK(clknet_leaf_62_clk),
    .D(net1688),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7801_ (.CLK(clknet_leaf_57_clk),
    .D(net1310),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7802_ (.CLK(clknet_leaf_40_clk),
    .D(net1745),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7803_ (.CLK(clknet_leaf_62_clk),
    .D(net1819),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7804_ (.CLK(clknet_leaf_37_clk),
    .D(net1095),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7805_ (.CLK(clknet_leaf_69_clk),
    .D(net1298),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7806_ (.CLK(clknet_leaf_59_clk),
    .D(net1231),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7807_ (.CLK(clknet_leaf_50_clk),
    .D(net1390),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7808_ (.CLK(clknet_leaf_71_clk),
    .D(net1370),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7809_ (.CLK(clknet_leaf_69_clk),
    .D(net989),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7810_ (.CLK(clknet_leaf_71_clk),
    .D(net1454),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7811_ (.CLK(clknet_leaf_54_clk),
    .D(net1520),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7812_ (.CLK(clknet_leaf_37_clk),
    .D(net1181),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7813_ (.CLK(clknet_leaf_35_clk),
    .D(net1721),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7814_ (.CLK(clknet_leaf_35_clk),
    .D(net1023),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7815_ (.CLK(clknet_leaf_35_clk),
    .D(net1414),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7816_ (.CLK(clknet_leaf_29_clk),
    .D(net1680),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7817_ (.CLK(clknet_leaf_20_clk),
    .D(net1684),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7818_ (.CLK(clknet_leaf_44_clk),
    .D(net1678),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7819_ (.CLK(clknet_leaf_68_clk),
    .D(net1430),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7820_ (.CLK(clknet_leaf_66_clk),
    .D(net1368),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7821_ (.CLK(clknet_leaf_41_clk),
    .D(net1548),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7822_ (.CLK(clknet_leaf_65_clk),
    .D(net1480),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7823_ (.CLK(clknet_leaf_71_clk),
    .D(net1388),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7824_ (.CLK(clknet_leaf_46_clk),
    .D(net1392),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7825_ (.CLK(clknet_leaf_41_clk),
    .D(net1554),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7826_ (.CLK(clknet_leaf_23_clk),
    .D(net1438),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7827_ (.CLK(clknet_leaf_25_clk),
    .D(net1494),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7828_ (.CLK(clknet_leaf_51_clk),
    .D(net1704),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7829_ (.CLK(clknet_leaf_44_clk),
    .D(net1795),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7830_ (.CLK(clknet_leaf_22_clk),
    .D(net987),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7831_ (.CLK(clknet_leaf_32_clk),
    .D(net1215),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7832_ (.CLK(clknet_leaf_59_clk),
    .D(net1588),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7833_ (.CLK(clknet_leaf_57_clk),
    .D(net1057),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7834_ (.CLK(clknet_leaf_40_clk),
    .D(net1492),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7835_ (.CLK(clknet_leaf_62_clk),
    .D(net1825),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7836_ (.CLK(clknet_leaf_40_clk),
    .D(net1648),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7837_ (.CLK(clknet_leaf_62_clk),
    .D(net1741),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7838_ (.CLK(clknet_leaf_57_clk),
    .D(net1225),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7839_ (.CLK(clknet_leaf_51_clk),
    .D(net1658),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7840_ (.CLK(clknet_leaf_70_clk),
    .D(net1692),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7841_ (.CLK(clknet_leaf_61_clk),
    .D(net1682),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7842_ (.CLK(clknet_leaf_70_clk),
    .D(net1396),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7843_ (.CLK(clknet_leaf_54_clk),
    .D(net1650),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7844_ (.CLK(clknet_leaf_6_clk),
    .D(_0604_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_src_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7845_ (.CLK(clknet_leaf_6_clk),
    .D(_0605_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7846_ (.CLK(clknet_leaf_4_clk),
    .D(_0606_),
    .Q(\U_DATAPATH.U_EX_MEM.i_mem_write_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7847_ (.CLK(clknet_leaf_4_clk),
    .D(_0607_),
    .Q(\U_DATAPATH.U_EX_MEM.i_result_src_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7848_ (.CLK(clknet_leaf_25_clk),
    .D(_0608_),
    .Q(\U_DATAPATH.U_EX_MEM.i_reg_write_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7849_ (.CLK(clknet_leaf_34_clk),
    .D(net802),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7850_ (.CLK(clknet_leaf_16_clk),
    .D(net947),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7851_ (.CLK(clknet_leaf_19_clk),
    .D(net993),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7852_ (.CLK(clknet_leaf_13_clk),
    .D(net895),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7853_ (.CLK(clknet_leaf_44_clk),
    .D(net2000),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7854_ (.CLK(clknet_leaf_9_clk),
    .D(net945),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7855_ (.CLK(clknet_leaf_13_clk),
    .D(net897),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7856_ (.CLK(clknet_leaf_9_clk),
    .D(net933),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7857_ (.CLK(clknet_leaf_3_clk),
    .D(net903),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7858_ (.CLK(clknet_leaf_4_clk),
    .D(net869),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7859_ (.CLK(clknet_leaf_3_clk),
    .D(net923),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7860_ (.CLK(clknet_leaf_11_clk),
    .D(net975),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7861_ (.CLK(clknet_leaf_15_clk),
    .D(net961),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7862_ (.CLK(clknet_leaf_15_clk),
    .D(net965),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7863_ (.CLK(clknet_leaf_41_clk),
    .D(_0623_),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7864_ (.CLK(clknet_leaf_10_clk),
    .D(net1332),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7865_ (.CLK(clknet_leaf_22_clk),
    .D(net714),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7866_ (.CLK(clknet_leaf_27_clk),
    .D(net1316),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7867_ (.CLK(clknet_leaf_34_clk),
    .D(net907),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7868_ (.CLK(clknet_leaf_53_clk),
    .D(net1133),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7869_ (.CLK(clknet_leaf_49_clk),
    .D(net943),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7870_ (.CLK(clknet_leaf_53_clk),
    .D(net1087),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7871_ (.CLK(clknet_leaf_48_clk),
    .D(net871),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7872_ (.CLK(clknet_leaf_58_clk),
    .D(net1005),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7873_ (.CLK(clknet_leaf_54_clk),
    .D(net1077),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7874_ (.CLK(clknet_leaf_53_clk),
    .D(net1109),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7875_ (.CLK(clknet_leaf_74_clk),
    .D(net672),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7876_ (.CLK(clknet_leaf_0_clk),
    .D(net1029),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7877_ (.CLK(clknet_leaf_1_clk),
    .D(net1811),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7878_ (.CLK(clknet_leaf_53_clk),
    .D(net1021),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7879_ (.CLK(clknet_leaf_24_clk),
    .D(net1358),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7880_ (.CLK(clknet_leaf_24_clk),
    .D(net628),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7881_ (.CLK(clknet_leaf_28_clk),
    .D(net883),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7882_ (.CLK(clknet_leaf_11_clk),
    .D(net979),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7883_ (.CLK(clknet_leaf_8_clk),
    .D(net875),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7884_ (.CLK(clknet_leaf_12_clk),
    .D(net929),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7885_ (.CLK(clknet_leaf_4_clk),
    .D(net644),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7886_ (.CLK(clknet_leaf_8_clk),
    .D(net885),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7887_ (.CLK(clknet_leaf_6_clk),
    .D(net836),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7888_ (.CLK(clknet_leaf_4_clk),
    .D(net846),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7889_ (.CLK(clknet_leaf_11_clk),
    .D(net844),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7890_ (.CLK(clknet_leaf_10_clk),
    .D(net690),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7891_ (.CLK(clknet_leaf_10_clk),
    .D(net1035),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7892_ (.CLK(clknet_leaf_10_clk),
    .D(net626),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7893_ (.CLK(clknet_leaf_10_clk),
    .D(net702),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7894_ (.CLK(clknet_leaf_27_clk),
    .D(net1097),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7895_ (.CLK(clknet_leaf_21_clk),
    .D(net881),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7896_ (.CLK(clknet_leaf_29_clk),
    .D(net860),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7897_ (.CLK(clknet_leaf_59_clk),
    .D(net977),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7898_ (.CLK(clknet_leaf_49_clk),
    .D(net957),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7899_ (.CLK(clknet_leaf_44_clk),
    .D(net1027),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7900_ (.CLK(clknet_leaf_63_clk),
    .D(net913),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7901_ (.CLK(clknet_leaf_50_clk),
    .D(net1049),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7902_ (.CLK(clknet_leaf_58_clk),
    .D(net1141),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7903_ (.CLK(clknet_leaf_58_clk),
    .D(net1209),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7904_ (.CLK(clknet_leaf_48_clk),
    .D(net1211),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7905_ (.CLK(clknet_leaf_66_clk),
    .D(net927),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7906_ (.CLK(clknet_leaf_72_clk),
    .D(net818),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7907_ (.CLK(clknet_leaf_65_clk),
    .D(net1171),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7908_ (.CLK(clknet_leaf_49_clk),
    .D(net963),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7909_ (.CLK(clknet_leaf_24_clk),
    .D(_0669_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7910_ (.CLK(clknet_leaf_24_clk),
    .D(_0670_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7911_ (.CLK(clknet_leaf_24_clk),
    .D(_0671_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7912_ (.CLK(clknet_leaf_24_clk),
    .D(_0672_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7913_ (.CLK(clknet_leaf_34_clk),
    .D(_0673_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7914_ (.CLK(clknet_leaf_23_clk),
    .D(_0674_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7915_ (.CLK(clknet_leaf_23_clk),
    .D(_0675_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7916_ (.CLK(clknet_leaf_23_clk),
    .D(_0676_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7917_ (.CLK(clknet_leaf_37_clk),
    .D(_0677_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7918_ (.CLK(clknet_leaf_31_clk),
    .D(_0678_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7919_ (.CLK(clknet_leaf_31_clk),
    .D(_0679_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7920_ (.CLK(clknet_leaf_32_clk),
    .D(_0680_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7921_ (.CLK(clknet_leaf_27_clk),
    .D(_0681_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7922_ (.CLK(clknet_leaf_26_clk),
    .D(_0682_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7923_ (.CLK(clknet_leaf_43_clk),
    .D(_0683_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7924_ (.CLK(clknet_leaf_68_clk),
    .D(_0684_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7925_ (.CLK(clknet_leaf_65_clk),
    .D(_0685_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7926_ (.CLK(clknet_leaf_45_clk),
    .D(_0686_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7927_ (.CLK(clknet_leaf_6_clk),
    .D(_0687_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7928_ (.CLK(clknet_leaf_65_clk),
    .D(_0688_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7929_ (.CLK(clknet_leaf_46_clk),
    .D(_0689_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7930_ (.CLK(clknet_leaf_45_clk),
    .D(_0690_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7931_ (.CLK(clknet_leaf_24_clk),
    .D(_0691_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7932_ (.CLK(clknet_leaf_26_clk),
    .D(_0692_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7933_ (.CLK(clknet_leaf_50_clk),
    .D(_0693_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7934_ (.CLK(clknet_leaf_47_clk),
    .D(_0694_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7935_ (.CLK(clknet_leaf_25_clk),
    .D(_0695_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7936_ (.CLK(clknet_leaf_29_clk),
    .D(_0696_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7937_ (.CLK(clknet_leaf_58_clk),
    .D(_0697_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7938_ (.CLK(clknet_leaf_58_clk),
    .D(_0698_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7939_ (.CLK(clknet_leaf_37_clk),
    .D(_0699_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7940_ (.CLK(clknet_leaf_62_clk),
    .D(_0700_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7941_ (.CLK(clknet_leaf_46_clk),
    .D(_0701_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7942_ (.CLK(clknet_leaf_62_clk),
    .D(_0702_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7943_ (.CLK(clknet_leaf_58_clk),
    .D(_0703_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7944_ (.CLK(clknet_leaf_49_clk),
    .D(_0704_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7945_ (.CLK(clknet_leaf_66_clk),
    .D(_0705_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7946_ (.CLK(clknet_leaf_67_clk),
    .D(_0706_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7947_ (.CLK(clknet_leaf_66_clk),
    .D(_0707_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7948_ (.CLK(clknet_leaf_53_clk),
    .D(_0708_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[31] ));
 sky130_fd_sc_hd__dfxtp_2 _7949_ (.CLK(clknet_leaf_37_clk),
    .D(_0709_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7950_ (.CLK(clknet_leaf_36_clk),
    .D(_0710_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7951_ (.CLK(clknet_leaf_31_clk),
    .D(_0711_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7952_ (.CLK(clknet_leaf_24_clk),
    .D(_0712_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7953_ (.CLK(clknet_leaf_27_clk),
    .D(_0713_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7954_ (.CLK(clknet_leaf_25_clk),
    .D(_0714_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7955_ (.CLK(clknet_leaf_43_clk),
    .D(_0715_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ));
 sky130_fd_sc_hd__dfxtp_2 _7956_ (.CLK(clknet_leaf_68_clk),
    .D(_0716_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7957_ (.CLK(clknet_leaf_65_clk),
    .D(_0717_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7958_ (.CLK(clknet_leaf_44_clk),
    .D(_0718_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7959_ (.CLK(clknet_leaf_6_clk),
    .D(_0719_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7960_ (.CLK(clknet_leaf_65_clk),
    .D(_0720_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7961_ (.CLK(clknet_leaf_30_clk),
    .D(_0721_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7962_ (.CLK(clknet_leaf_45_clk),
    .D(_0722_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7963_ (.CLK(clknet_leaf_27_clk),
    .D(_0723_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7964_ (.CLK(clknet_leaf_26_clk),
    .D(_0724_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[15] ));
 sky130_fd_sc_hd__dfxtp_2 _7965_ (.CLK(clknet_leaf_48_clk),
    .D(_0725_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7966_ (.CLK(clknet_leaf_47_clk),
    .D(_0726_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7967_ (.CLK(clknet_leaf_25_clk),
    .D(_0727_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7968_ (.CLK(clknet_leaf_29_clk),
    .D(_0728_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7969_ (.CLK(clknet_leaf_58_clk),
    .D(_0729_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7970_ (.CLK(clknet_leaf_55_clk),
    .D(_0730_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[21] ));
 sky130_fd_sc_hd__dfxtp_2 _7971_ (.CLK(clknet_leaf_40_clk),
    .D(_0731_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7972_ (.CLK(clknet_leaf_63_clk),
    .D(_0732_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[23] ));
 sky130_fd_sc_hd__dfxtp_2 _7973_ (.CLK(clknet_leaf_46_clk),
    .D(_0733_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7974_ (.CLK(clknet_leaf_62_clk),
    .D(_0734_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7975_ (.CLK(clknet_leaf_58_clk),
    .D(_0735_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7976_ (.CLK(clknet_leaf_53_clk),
    .D(_0736_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7977_ (.CLK(clknet_leaf_66_clk),
    .D(_0737_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7978_ (.CLK(clknet_leaf_67_clk),
    .D(_0738_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7979_ (.CLK(clknet_leaf_66_clk),
    .D(_0739_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7980_ (.CLK(clknet_leaf_53_clk),
    .D(_0740_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7981_ (.CLK(clknet_leaf_22_clk),
    .D(_0741_),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7982_ (.CLK(clknet_leaf_22_clk),
    .D(_0742_),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7983_ (.CLK(clknet_leaf_23_clk),
    .D(_0743_),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7984_ (.CLK(clknet_leaf_22_clk),
    .D(_0744_),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7985_ (.CLK(clknet_leaf_6_clk),
    .D(_0745_),
    .Q(\U_DATAPATH.U_ID_EX.o_addr_src_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7986_ (.CLK(clknet_leaf_6_clk),
    .D(_0746_),
    .Q(\U_CONTROL_UNIT.i_branch_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7987_ (.CLK(clknet_leaf_6_clk),
    .D(_0747_),
    .Q(\U_CONTROL_UNIT.i_jump_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7988_ (.CLK(clknet_leaf_41_clk),
    .D(_0748_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7989_ (.CLK(clknet_leaf_44_clk),
    .D(net2152),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7990_ (.CLK(clknet_leaf_34_clk),
    .D(_0750_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7991_ (.CLK(clknet_leaf_16_clk),
    .D(_0751_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7992_ (.CLK(clknet_leaf_18_clk),
    .D(_0752_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7993_ (.CLK(clknet_leaf_11_clk),
    .D(_0753_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7994_ (.CLK(clknet_leaf_43_clk),
    .D(_0754_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7995_ (.CLK(clknet_leaf_8_clk),
    .D(_0755_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7996_ (.CLK(clknet_leaf_12_clk),
    .D(_0756_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7997_ (.CLK(clknet_leaf_28_clk),
    .D(_0757_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7998_ (.CLK(clknet_leaf_3_clk),
    .D(_0758_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7999_ (.CLK(clknet_leaf_4_clk),
    .D(_0759_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8000_ (.CLK(clknet_leaf_12_clk),
    .D(_0760_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8001_ (.CLK(clknet_leaf_9_clk),
    .D(_0761_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8002_ (.CLK(clknet_leaf_10_clk),
    .D(_0762_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8003_ (.CLK(clknet_leaf_15_clk),
    .D(_0763_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8004_ (.CLK(clknet_leaf_41_clk),
    .D(_0764_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8005_ (.CLK(clknet_leaf_10_clk),
    .D(_0765_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8006_ (.CLK(clknet_leaf_22_clk),
    .D(_0766_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8007_ (.CLK(clknet_leaf_27_clk),
    .D(_0767_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8008_ (.CLK(clknet_leaf_34_clk),
    .D(_0768_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8009_ (.CLK(clknet_leaf_53_clk),
    .D(_0769_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8010_ (.CLK(clknet_leaf_49_clk),
    .D(_0770_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8011_ (.CLK(clknet_leaf_53_clk),
    .D(_0771_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8012_ (.CLK(clknet_leaf_50_clk),
    .D(_0772_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8013_ (.CLK(clknet_leaf_58_clk),
    .D(_0773_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8014_ (.CLK(clknet_leaf_54_clk),
    .D(_0774_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8015_ (.CLK(clknet_leaf_53_clk),
    .D(_0775_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8016_ (.CLK(clknet_leaf_0_clk),
    .D(_0776_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8017_ (.CLK(clknet_leaf_0_clk),
    .D(_0777_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8018_ (.CLK(clknet_leaf_0_clk),
    .D(_0778_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8019_ (.CLK(clknet_leaf_53_clk),
    .D(_0779_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8020_ (.CLK(clknet_leaf_23_clk),
    .D(net686),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8021_ (.CLK(clknet_leaf_23_clk),
    .D(net682),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8022_ (.CLK(clknet_leaf_23_clk),
    .D(_0782_),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8023_ (.CLK(clknet_leaf_23_clk),
    .D(net674),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8024_ (.CLK(clknet_leaf_34_clk),
    .D(net734),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8025_ (.CLK(clknet_leaf_16_clk),
    .D(net776),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8026_ (.CLK(clknet_leaf_18_clk),
    .D(net754),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8027_ (.CLK(clknet_leaf_11_clk),
    .D(net638),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8028_ (.CLK(clknet_leaf_43_clk),
    .D(net854),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8029_ (.CLK(clknet_leaf_8_clk),
    .D(net694),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8030_ (.CLK(clknet_leaf_12_clk),
    .D(net642),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8031_ (.CLK(clknet_leaf_8_clk),
    .D(net750),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8032_ (.CLK(clknet_leaf_3_clk),
    .D(net762),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8033_ (.CLK(clknet_leaf_4_clk),
    .D(net804),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8034_ (.CLK(clknet_leaf_3_clk),
    .D(net748),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8035_ (.CLK(clknet_leaf_9_clk),
    .D(net664),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8036_ (.CLK(clknet_leaf_11_clk),
    .D(net668),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8037_ (.CLK(clknet_leaf_16_clk),
    .D(net650),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8038_ (.CLK(clknet_leaf_41_clk),
    .D(net756),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8039_ (.CLK(clknet_leaf_10_clk),
    .D(net812),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8040_ (.CLK(clknet_leaf_22_clk),
    .D(net728),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8041_ (.CLK(clknet_leaf_27_clk),
    .D(net822),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8042_ (.CLK(clknet_leaf_34_clk),
    .D(net770),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8043_ (.CLK(clknet_leaf_53_clk),
    .D(net794),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8044_ (.CLK(clknet_leaf_49_clk),
    .D(net764),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8045_ (.CLK(clknet_leaf_53_clk),
    .D(net774),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8046_ (.CLK(clknet_leaf_48_clk),
    .D(net744),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8047_ (.CLK(clknet_leaf_58_clk),
    .D(net808),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8048_ (.CLK(clknet_leaf_55_clk),
    .D(net658),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8049_ (.CLK(clknet_leaf_53_clk),
    .D(net887),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8050_ (.CLK(clknet_leaf_0_clk),
    .D(net634),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8051_ (.CLK(clknet_leaf_0_clk),
    .D(net824),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8052_ (.CLK(clknet_leaf_1_clk),
    .D(net700),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8053_ (.CLK(clknet_leaf_53_clk),
    .D(net792),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8054_ (.CLK(clknet_leaf_29_clk),
    .D(net2356),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8055_ (.CLK(clknet_leaf_47_clk),
    .D(_0815_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8056_ (.CLK(clknet_leaf_32_clk),
    .D(net2335),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8057_ (.CLK(clknet_leaf_32_clk),
    .D(_0817_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8058_ (.CLK(clknet_leaf_27_clk),
    .D(net2372),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8059_ (.CLK(clknet_leaf_27_clk),
    .D(net2322),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8060_ (.CLK(clknet_leaf_7_clk),
    .D(net2332),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8061_ (.CLK(clknet_leaf_68_clk),
    .D(_0821_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8062_ (.CLK(clknet_leaf_65_clk),
    .D(_0822_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8063_ (.CLK(clknet_leaf_28_clk),
    .D(net2348),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8064_ (.CLK(clknet_leaf_65_clk),
    .D(net2340),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8065_ (.CLK(clknet_leaf_65_clk),
    .D(_0825_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8066_ (.CLK(clknet_leaf_28_clk),
    .D(_0826_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8067_ (.CLK(clknet_leaf_29_clk),
    .D(_0827_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8068_ (.CLK(clknet_leaf_27_clk),
    .D(_0828_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8069_ (.CLK(clknet_leaf_26_clk),
    .D(_0829_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8070_ (.CLK(clknet_leaf_48_clk),
    .D(_0830_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8071_ (.CLK(clknet_leaf_47_clk),
    .D(net2325),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8072_ (.CLK(clknet_leaf_27_clk),
    .D(net2338),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8073_ (.CLK(clknet_leaf_30_clk),
    .D(net2368),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8074_ (.CLK(clknet_leaf_63_clk),
    .D(_0834_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8075_ (.CLK(clknet_leaf_63_clk),
    .D(net2342),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8076_ (.CLK(clknet_leaf_47_clk),
    .D(_0836_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8077_ (.CLK(clknet_leaf_62_clk),
    .D(net2312),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8078_ (.CLK(clknet_leaf_48_clk),
    .D(_0838_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8079_ (.CLK(clknet_leaf_62_clk),
    .D(_0839_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8080_ (.CLK(clknet_leaf_63_clk),
    .D(net2352),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8081_ (.CLK(clknet_leaf_48_clk),
    .D(net2329),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8082_ (.CLK(clknet_leaf_67_clk),
    .D(_0842_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8083_ (.CLK(clknet_leaf_67_clk),
    .D(_0843_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8084_ (.CLK(clknet_leaf_65_clk),
    .D(_0844_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8085_ (.CLK(clknet_3_3_0_clk),
    .D(_0845_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8086_ (.CLK(clknet_leaf_51_clk),
    .D(_0846_),
    .Q(\U_DATAPATH.U_EX_MEM.o_result_src_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8087_ (.CLK(clknet_leaf_12_clk),
    .D(net1436),
    .Q(\U_DATAPATH.U_EX_MEM.o_result_src_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8088_ (.CLK(clknet_leaf_22_clk),
    .D(net1940),
    .Q(\U_DATAPATH.U_EX_MEM.o_reg_write_M ));
 sky130_fd_sc_hd__dfxtp_1 _8089_ (.CLK(clknet_leaf_55_clk),
    .D(_0849_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8090_ (.CLK(clknet_leaf_2_clk),
    .D(_0850_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8091_ (.CLK(clknet_leaf_2_clk),
    .D(_0851_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8092_ (.CLK(clknet_leaf_35_clk),
    .D(_0852_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8093_ (.CLK(clknet_leaf_34_clk),
    .D(_0853_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8094_ (.CLK(clknet_leaf_17_clk),
    .D(_0854_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8095_ (.CLK(clknet_leaf_14_clk),
    .D(_0855_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8096_ (.CLK(clknet_leaf_56_clk),
    .D(_0856_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8097_ (.CLK(clknet_leaf_0_clk),
    .D(_0857_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8098_ (.CLK(clknet_leaf_15_clk),
    .D(_0858_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8099_ (.CLK(clknet_leaf_35_clk),
    .D(_0859_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8100_ (.CLK(clknet_leaf_74_clk),
    .D(_0860_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8101_ (.CLK(clknet_leaf_15_clk),
    .D(_0861_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8102_ (.CLK(clknet_leaf_57_clk),
    .D(_0862_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8103_ (.CLK(clknet_leaf_14_clk),
    .D(_0863_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8104_ (.CLK(clknet_leaf_15_clk),
    .D(_0864_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8105_ (.CLK(clknet_leaf_13_clk),
    .D(_0865_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8106_ (.CLK(clknet_leaf_14_clk),
    .D(net2156),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8107_ (.CLK(clknet_leaf_21_clk),
    .D(_0867_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8108_ (.CLK(clknet_leaf_14_clk),
    .D(_0868_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8109_ (.CLK(clknet_leaf_74_clk),
    .D(_0869_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8110_ (.CLK(clknet_leaf_74_clk),
    .D(_0870_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8111_ (.CLK(clknet_leaf_18_clk),
    .D(_0871_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8112_ (.CLK(clknet_leaf_61_clk),
    .D(_0872_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8113_ (.CLK(clknet_leaf_38_clk),
    .D(_0873_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8114_ (.CLK(clknet_leaf_52_clk),
    .D(_0874_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8115_ (.CLK(clknet_leaf_74_clk),
    .D(_0875_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8116_ (.CLK(clknet_leaf_42_clk),
    .D(_0876_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8117_ (.CLK(clknet_leaf_74_clk),
    .D(_0877_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8118_ (.CLK(clknet_leaf_70_clk),
    .D(_0878_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[29] ));
 sky130_fd_sc_hd__dfxtp_2 _8119_ (.CLK(clknet_leaf_53_clk),
    .D(_0879_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8120_ (.CLK(clknet_leaf_60_clk),
    .D(_0880_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8121_ (.CLK(clknet_leaf_3_clk),
    .D(net842),
    .Q(\U_DATAPATH.U_EX_MEM.o_mem_write_M ));
 sky130_fd_sc_hd__dfxtp_1 _8122_ (.CLK(clknet_leaf_22_clk),
    .D(net740),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _8123_ (.CLK(clknet_leaf_35_clk),
    .D(net622),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_2 _8124_ (.CLK(clknet_leaf_1_clk),
    .D(net850),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _8125_ (.CLK(clknet_leaf_23_clk),
    .D(net732),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ));
 sky130_fd_sc_hd__dfxtp_4 _8126_ (.CLK(clknet_leaf_33_clk),
    .D(net2119),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ));
 sky130_fd_sc_hd__dfxtp_4 _8127_ (.CLK(clknet_leaf_33_clk),
    .D(net2040),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ));
 sky130_fd_sc_hd__dfxtp_4 _8128_ (.CLK(clknet_leaf_33_clk),
    .D(net2101),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ));
 sky130_fd_sc_hd__dfxtp_4 _8129_ (.CLK(clknet_leaf_33_clk),
    .D(net2113),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8130_ (.CLK(clknet_leaf_34_clk),
    .D(net742),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8131_ (.CLK(clknet_leaf_16_clk),
    .D(net752),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8132_ (.CLK(clknet_leaf_18_clk),
    .D(net724),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8133_ (.CLK(clknet_leaf_11_clk),
    .D(net738),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8134_ (.CLK(clknet_leaf_43_clk),
    .D(net826),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8135_ (.CLK(clknet_leaf_8_clk),
    .D(net746),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8136_ (.CLK(clknet_leaf_12_clk),
    .D(net718),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8137_ (.CLK(clknet_leaf_28_clk),
    .D(net688),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8138_ (.CLK(clknet_leaf_4_clk),
    .D(net660),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8139_ (.CLK(clknet_leaf_4_clk),
    .D(net758),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8140_ (.CLK(clknet_leaf_12_clk),
    .D(net620),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8141_ (.CLK(clknet_leaf_9_clk),
    .D(net782),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8142_ (.CLK(clknet_leaf_10_clk),
    .D(net630),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8143_ (.CLK(clknet_leaf_16_clk),
    .D(net780),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8144_ (.CLK(clknet_leaf_42_clk),
    .D(net696),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8145_ (.CLK(clknet_leaf_10_clk),
    .D(net786),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8146_ (.CLK(clknet_leaf_22_clk),
    .D(net712),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8147_ (.CLK(clknet_leaf_27_clk),
    .D(net810),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8148_ (.CLK(clknet_leaf_34_clk),
    .D(net766),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8149_ (.CLK(clknet_leaf_52_clk),
    .D(net692),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8150_ (.CLK(clknet_leaf_53_clk),
    .D(net636),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8151_ (.CLK(clknet_leaf_52_clk),
    .D(net684),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8152_ (.CLK(clknet_leaf_50_clk),
    .D(net654),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8153_ (.CLK(clknet_leaf_54_clk),
    .D(net830),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8154_ (.CLK(clknet_leaf_55_clk),
    .D(net778),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8155_ (.CLK(clknet_leaf_53_clk),
    .D(net840),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8156_ (.CLK(clknet_leaf_72_clk),
    .D(net646),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8157_ (.CLK(clknet_leaf_0_clk),
    .D(net806),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8158_ (.CLK(clknet_leaf_1_clk),
    .D(net708),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8159_ (.CLK(clknet_leaf_52_clk),
    .D(net698),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8160_ (.CLK(clknet_leaf_41_clk),
    .D(net796),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8161_ (.CLK(clknet_leaf_42_clk),
    .D(net800),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8162_ (.CLK(clknet_leaf_34_clk),
    .D(net772),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8163_ (.CLK(clknet_leaf_16_clk),
    .D(net798),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8164_ (.CLK(clknet_leaf_18_clk),
    .D(net730),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8165_ (.CLK(clknet_leaf_11_clk),
    .D(net760),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8166_ (.CLK(clknet_leaf_43_clk),
    .D(net784),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8167_ (.CLK(clknet_leaf_7_clk),
    .D(net706),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8168_ (.CLK(clknet_leaf_12_clk),
    .D(net710),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8169_ (.CLK(clknet_leaf_28_clk),
    .D(net828),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8170_ (.CLK(clknet_leaf_4_clk),
    .D(net666),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8171_ (.CLK(clknet_leaf_5_clk),
    .D(net670),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8172_ (.CLK(clknet_leaf_12_clk),
    .D(net704),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8173_ (.CLK(clknet_leaf_7_clk),
    .D(net834),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8174_ (.CLK(clknet_leaf_11_clk),
    .D(net820),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8175_ (.CLK(clknet_leaf_10_clk),
    .D(net632),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8176_ (.CLK(clknet_leaf_42_clk),
    .D(net720),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8177_ (.CLK(clknet_leaf_10_clk),
    .D(net832),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8178_ (.CLK(clknet_leaf_22_clk),
    .D(net722),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8179_ (.CLK(clknet_leaf_27_clk),
    .D(net788),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8180_ (.CLK(clknet_leaf_35_clk),
    .D(net648),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8181_ (.CLK(clknet_leaf_53_clk),
    .D(net814),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8182_ (.CLK(clknet_leaf_49_clk),
    .D(net726),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8183_ (.CLK(clknet_leaf_52_clk),
    .D(net678),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8184_ (.CLK(clknet_leaf_47_clk),
    .D(net652),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8185_ (.CLK(clknet_leaf_54_clk),
    .D(net816),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8186_ (.CLK(clknet_leaf_55_clk),
    .D(net640),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8187_ (.CLK(clknet_leaf_52_clk),
    .D(net848),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8188_ (.CLK(clknet_leaf_72_clk),
    .D(net656),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8189_ (.CLK(clknet_leaf_0_clk),
    .D(net838),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8190_ (.CLK(clknet_leaf_5_clk),
    .D(net676),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8191_ (.CLK(clknet_leaf_52_clk),
    .D(net680),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8192_ (.CLK(clknet_leaf_42_clk),
    .D(_0952_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8193_ (.CLK(clknet_leaf_51_clk),
    .D(_0953_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8194_ (.CLK(clknet_leaf_35_clk),
    .D(_0954_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8195_ (.CLK(clknet_leaf_19_clk),
    .D(_0955_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8196_ (.CLK(clknet_leaf_18_clk),
    .D(_0956_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8197_ (.CLK(clknet_leaf_14_clk),
    .D(_0957_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8198_ (.CLK(clknet_leaf_43_clk),
    .D(_0958_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[6] ));
 sky130_fd_sc_hd__dfxtp_2 _8199_ (.CLK(clknet_leaf_23_clk),
    .D(_0959_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8200_ (.CLK(clknet_leaf_13_clk),
    .D(_0960_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[8] ));
 sky130_fd_sc_hd__dfxtp_2 _8201_ (.CLK(clknet_leaf_34_clk),
    .D(_0961_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8202_ (.CLK(clknet_leaf_1_clk),
    .D(_0962_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8203_ (.CLK(clknet_leaf_73_clk),
    .D(_0963_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8204_ (.CLK(clknet_leaf_14_clk),
    .D(_0964_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8205_ (.CLK(clknet_leaf_43_clk),
    .D(_0965_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8206_ (.CLK(clknet_leaf_4_clk),
    .D(_0966_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[14] ));
 sky130_fd_sc_hd__dfxtp_2 _8207_ (.CLK(clknet_leaf_0_clk),
    .D(_0967_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8208_ (.CLK(clknet_leaf_43_clk),
    .D(_0968_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8209_ (.CLK(clknet_leaf_17_clk),
    .D(_0969_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8210_ (.CLK(clknet_leaf_39_clk),
    .D(_0970_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[18] ));
 sky130_fd_sc_hd__dfxtp_4 _8211_ (.CLK(clknet_leaf_73_clk),
    .D(_0971_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8212_ (.CLK(clknet_leaf_39_clk),
    .D(_0972_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8213_ (.CLK(clknet_leaf_42_clk),
    .D(_0973_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8214_ (.CLK(clknet_leaf_2_clk),
    .D(_0974_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8215_ (.CLK(clknet_leaf_52_clk),
    .D(_0975_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[23] ));
 sky130_fd_sc_hd__dfxtp_2 _8216_ (.CLK(clknet_leaf_17_clk),
    .D(_0976_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8217_ (.CLK(clknet_leaf_56_clk),
    .D(_0977_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8218_ (.CLK(clknet_leaf_55_clk),
    .D(_0978_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8219_ (.CLK(clknet_leaf_52_clk),
    .D(_0979_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8220_ (.CLK(clknet_leaf_74_clk),
    .D(_0980_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8221_ (.CLK(clknet_leaf_1_clk),
    .D(_0981_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8222_ (.CLK(clknet_leaf_1_clk),
    .D(_0982_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8223_ (.CLK(clknet_leaf_56_clk),
    .D(_0983_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8224_ (.CLK(net521),
    .D(_0984_),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_1 _8225_ (.CLK(net522),
    .D(_0985_),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_2 _8226_ (.CLK(net523),
    .D(_0986_),
    .Q(net152));
 sky130_fd_sc_hd__dfxtp_1 _8227_ (.CLK(net524),
    .D(_0987_),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_1 _8228_ (.CLK(net525),
    .D(_0988_),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_1 _8229_ (.CLK(net526),
    .D(_0989_),
    .Q(net157));
 sky130_fd_sc_hd__dfxtp_2 _8230_ (.CLK(net527),
    .D(_0990_),
    .Q(net158));
 sky130_fd_sc_hd__dfxtp_1 _8231_ (.CLK(net528),
    .D(_0991_),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_1 _8232_ (.CLK(net529),
    .D(_0992_),
    .Q(net160));
 sky130_fd_sc_hd__dfxtp_1 _8233_ (.CLK(net530),
    .D(_0993_),
    .Q(net161));
 sky130_fd_sc_hd__dfxtp_1 _8234_ (.CLK(net531),
    .D(_0994_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_1 _8235_ (.CLK(net532),
    .D(_0995_),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_1 _8236_ (.CLK(net533),
    .D(_0996_),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_1 _8237_ (.CLK(net534),
    .D(_0997_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_4 _8238_ (.CLK(net535),
    .D(_0998_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_4 _8239_ (.CLK(net536),
    .D(_0999_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_2 _8240_ (.CLK(net537),
    .D(_1000_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_2 _8241_ (.CLK(net538),
    .D(_1001_),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_1 _8242_ (.CLK(net539),
    .D(_1002_),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_1 _8243_ (.CLK(net540),
    .D(_1003_),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_2 _8244_ (.CLK(net541),
    .D(_1004_),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_1 _8245_ (.CLK(net542),
    .D(_1005_),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_1 _8246_ (.CLK(net543),
    .D(_1006_),
    .Q(net144));
 sky130_fd_sc_hd__dfxtp_1 _8247_ (.CLK(net544),
    .D(_1007_),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_1 _8248_ (.CLK(net545),
    .D(_1008_),
    .Q(net146));
 sky130_fd_sc_hd__dfxtp_1 _8249_ (.CLK(net546),
    .D(_1009_),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_2 _8250_ (.CLK(net547),
    .D(_1010_),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_1 _8251_ (.CLK(net548),
    .D(_1011_),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_1 _8252_ (.CLK(net549),
    .D(_1012_),
    .Q(net150));
 sky130_fd_sc_hd__dfxtp_1 _8253_ (.CLK(net550),
    .D(_1013_),
    .Q(net151));
 sky130_fd_sc_hd__dfxtp_1 _8254_ (.CLK(net551),
    .D(_1014_),
    .Q(net153));
 sky130_fd_sc_hd__dfxtp_1 _8255_ (.CLK(net552),
    .D(_1015_),
    .Q(net154));
 sky130_fd_sc_hd__dfxtp_1 _8256_ (.CLK(clknet_leaf_42_clk),
    .D(_0069_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8257_ (.CLK(clknet_leaf_42_clk),
    .D(_0080_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8258_ (.CLK(clknet_leaf_31_clk),
    .D(net1781),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8259_ (.CLK(clknet_leaf_16_clk),
    .D(_0094_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8260_ (.CLK(clknet_leaf_10_clk),
    .D(_0095_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8261_ (.CLK(clknet_leaf_26_clk),
    .D(_0096_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8262_ (.CLK(clknet_leaf_51_clk),
    .D(_0097_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8263_ (.CLK(clknet_leaf_68_clk),
    .D(_0098_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8264_ (.CLK(clknet_leaf_5_clk),
    .D(_0099_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8265_ (.CLK(clknet_leaf_28_clk),
    .D(net1920),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8266_ (.CLK(clknet_leaf_4_clk),
    .D(_0070_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8267_ (.CLK(clknet_leaf_5_clk),
    .D(_0071_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8268_ (.CLK(clknet_leaf_47_clk),
    .D(net1823),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8269_ (.CLK(clknet_leaf_45_clk),
    .D(_0073_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8270_ (.CLK(clknet_leaf_27_clk),
    .D(_0074_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8271_ (.CLK(clknet_leaf_16_clk),
    .D(_0075_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8272_ (.CLK(clknet_leaf_51_clk),
    .D(_0076_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8273_ (.CLK(clknet_leaf_48_clk),
    .D(_0077_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8274_ (.CLK(clknet_leaf_25_clk),
    .D(_0078_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8275_ (.CLK(clknet_leaf_27_clk),
    .D(net768),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8276_ (.CLK(clknet_leaf_63_clk),
    .D(_0081_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8277_ (.CLK(clknet_leaf_55_clk),
    .D(_0082_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8278_ (.CLK(clknet_leaf_40_clk),
    .D(_0083_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8279_ (.CLK(clknet_leaf_62_clk),
    .D(_0084_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8280_ (.CLK(clknet_leaf_47_clk),
    .D(_0085_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8281_ (.CLK(clknet_leaf_62_clk),
    .D(_0086_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8282_ (.CLK(clknet_leaf_55_clk),
    .D(_0087_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8283_ (.CLK(clknet_leaf_52_clk),
    .D(_0088_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8284_ (.CLK(clknet_leaf_0_clk),
    .D(_0089_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8285_ (.CLK(clknet_leaf_67_clk),
    .D(_0090_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8286_ (.CLK(clknet_leaf_0_clk),
    .D(_0092_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8287_ (.CLK(clknet_leaf_52_clk),
    .D(net624),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[31] ));
 sky130_fd_sc_hd__dfxtp_2 _8288_ (.CLK(net553),
    .D(_1016_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_1 _8289_ (.CLK(clknet_leaf_22_clk),
    .D(_1017_),
    .Q(\U_DATAPATH.U_EX_MEM.i_funct3_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8290_ (.CLK(clknet_leaf_21_clk),
    .D(_1018_),
    .Q(\U_DATAPATH.U_EX_MEM.i_funct3_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8291_ (.CLK(clknet_leaf_3_clk),
    .D(_1019_),
    .Q(\U_DATAPATH.U_EX_MEM.i_funct3_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8292_ (.CLK(net554),
    .D(_0069_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_2 _8293_ (.CLK(net555),
    .D(_0080_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_4 _8294_ (.CLK(net556),
    .D(_0091_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_2 _8295_ (.CLK(net557),
    .D(_0094_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_2 _8296_ (.CLK(net558),
    .D(_0095_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_2 _8297_ (.CLK(net559),
    .D(_0096_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_2 _8298_ (.CLK(net560),
    .D(_0097_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_2 _8299_ (.CLK(net561),
    .D(_0098_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_2 _8300_ (.CLK(net562),
    .D(_0099_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_2 _8301_ (.CLK(net563),
    .D(_0100_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_2 _8302_ (.CLK(net564),
    .D(_0070_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_2 _8303_ (.CLK(net565),
    .D(_0071_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_4 _8304_ (.CLK(net566),
    .D(_0072_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_2 _8305_ (.CLK(net567),
    .D(_0073_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_2 _8306_ (.CLK(net568),
    .D(_0074_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_2 _8307_ (.CLK(net569),
    .D(_0075_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_2 _8308_ (.CLK(net570),
    .D(_0076_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_2 _8309_ (.CLK(net571),
    .D(_0077_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_2 _8310_ (.CLK(net572),
    .D(_0078_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_2 _8311_ (.CLK(net573),
    .D(_0079_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _8312_ (.CLK(net574),
    .D(_0081_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_2 _8313_ (.CLK(net575),
    .D(_0082_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _8314_ (.CLK(net576),
    .D(_0083_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_2 _8315_ (.CLK(net577),
    .D(_0084_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_4 _8316_ (.CLK(net578),
    .D(_0085_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_2 _8317_ (.CLK(net579),
    .D(_0086_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _8318_ (.CLK(net580),
    .D(_0087_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _8319_ (.CLK(net581),
    .D(_0088_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_4 _8320_ (.CLK(net582),
    .D(_0089_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_4 _8321_ (.CLK(net583),
    .D(_0090_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_1 _8322_ (.CLK(net584),
    .D(_0092_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_2 _8323_ (.CLK(net585),
    .D(_0093_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _8324_ (.CLK(net586),
    .D(_0032_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8325_ (.CLK(net587),
    .D(_0043_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8326_ (.CLK(net588),
    .D(_0054_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8327_ (.CLK(net589),
    .D(_0057_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8328_ (.CLK(net590),
    .D(_0058_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8329_ (.CLK(net591),
    .D(_0059_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8330_ (.CLK(net592),
    .D(_0060_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8331_ (.CLK(net593),
    .D(_0061_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8332_ (.CLK(net594),
    .D(_0062_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8333_ (.CLK(net595),
    .D(_0063_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8334_ (.CLK(net596),
    .D(_0033_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8335_ (.CLK(net597),
    .D(_0034_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8336_ (.CLK(net598),
    .D(_0035_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8337_ (.CLK(net599),
    .D(_0036_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8338_ (.CLK(net600),
    .D(_0037_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8339_ (.CLK(net601),
    .D(_0038_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8340_ (.CLK(net602),
    .D(_0039_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8341_ (.CLK(net603),
    .D(_0040_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8342_ (.CLK(net604),
    .D(_0041_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8343_ (.CLK(net605),
    .D(_0042_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8344_ (.CLK(net606),
    .D(_0044_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8345_ (.CLK(net607),
    .D(_0045_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8346_ (.CLK(net608),
    .D(_0046_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8347_ (.CLK(net609),
    .D(_0047_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8348_ (.CLK(net610),
    .D(_0048_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8349_ (.CLK(net611),
    .D(_0049_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8350_ (.CLK(net612),
    .D(_0050_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8351_ (.CLK(net613),
    .D(_0051_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8352_ (.CLK(net614),
    .D(_0052_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8353_ (.CLK(net615),
    .D(_0053_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8354_ (.CLK(net616),
    .D(_0055_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8355_ (.CLK(net617),
    .D(_0056_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8356_ (.CLK(clknet_leaf_38_clk),
    .D(net925),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8357_ (.CLK(clknet_leaf_39_clk),
    .D(net858),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8358_ (.CLK(clknet_leaf_38_clk),
    .D(net1558),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8359_ (.CLK(clknet_leaf_33_clk),
    .D(net1107),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8360_ (.CLK(clknet_leaf_29_clk),
    .D(net1526),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8361_ (.CLK(clknet_leaf_19_clk),
    .D(net1638),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8362_ (.CLK(clknet_leaf_43_clk),
    .D(net919),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8363_ (.CLK(clknet_leaf_68_clk),
    .D(net1115),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8364_ (.CLK(clknet_leaf_5_clk),
    .D(net1340),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8365_ (.CLK(clknet_leaf_45_clk),
    .D(net1165),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8366_ (.CLK(clknet_leaf_4_clk),
    .D(net1197),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8367_ (.CLK(clknet_leaf_72_clk),
    .D(net1067),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8368_ (.CLK(clknet_leaf_46_clk),
    .D(net1460),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8369_ (.CLK(clknet_leaf_41_clk),
    .D(net1386),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8370_ (.CLK(clknet_leaf_25_clk),
    .D(net1376),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8371_ (.CLK(clknet_leaf_16_clk),
    .D(net1153),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8372_ (.CLK(clknet_leaf_52_clk),
    .D(net1540),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8373_ (.CLK(clknet_leaf_48_clk),
    .D(net1328),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8374_ (.CLK(clknet_leaf_20_clk),
    .D(net953),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8375_ (.CLK(clknet_leaf_27_clk),
    .D(net1348),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8376_ (.CLK(clknet_leaf_60_clk),
    .D(net1099),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8377_ (.CLK(clknet_leaf_56_clk),
    .D(net1277),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8378_ (.CLK(clknet_leaf_40_clk),
    .D(net1233),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8379_ (.CLK(clknet_leaf_61_clk),
    .D(net1516),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8380_ (.CLK(clknet_leaf_31_clk),
    .D(net1729),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8381_ (.CLK(clknet_leaf_69_clk),
    .D(net1045),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8382_ (.CLK(clknet_leaf_59_clk),
    .D(net1039),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8383_ (.CLK(clknet_leaf_51_clk),
    .D(net1590),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8384_ (.CLK(clknet_leaf_72_clk),
    .D(net1059),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8385_ (.CLK(clknet_leaf_70_clk),
    .D(net1344),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8386_ (.CLK(clknet_leaf_70_clk),
    .D(net1426),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8387_ (.CLK(clknet_leaf_55_clk),
    .D(net1594),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8388_ (.CLK(clknet_leaf_37_clk),
    .D(net1873),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8389_ (.CLK(clknet_leaf_39_clk),
    .D(net1769),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8390_ (.CLK(clknet_leaf_37_clk),
    .D(net2137),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8391_ (.CLK(clknet_leaf_32_clk),
    .D(net1773),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8392_ (.CLK(clknet_leaf_31_clk),
    .D(net1891),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8393_ (.CLK(clknet_leaf_19_clk),
    .D(net1902),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8394_ (.CLK(clknet_leaf_43_clk),
    .D(net1676),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8395_ (.CLK(clknet_leaf_62_clk),
    .D(net1973),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8396_ (.CLK(clknet_leaf_66_clk),
    .D(net1975),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8397_ (.CLK(clknet_leaf_42_clk),
    .D(net1954),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8398_ (.CLK(clknet_leaf_5_clk),
    .D(net1956),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8399_ (.CLK(clknet_leaf_71_clk),
    .D(net1881),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8400_ (.CLK(clknet_leaf_46_clk),
    .D(net1711),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8401_ (.CLK(clknet_leaf_41_clk),
    .D(net1990),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8402_ (.CLK(clknet_leaf_20_clk),
    .D(net1596),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8403_ (.CLK(clknet_leaf_16_clk),
    .D(net1926),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8404_ (.CLK(clknet_leaf_52_clk),
    .D(net1987),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8405_ (.CLK(clknet_leaf_44_clk),
    .D(net1885),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8406_ (.CLK(clknet_leaf_20_clk),
    .D(net1777),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8407_ (.CLK(clknet_leaf_29_clk),
    .D(net1942),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8408_ (.CLK(clknet_leaf_60_clk),
    .D(net1686),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8409_ (.CLK(clknet_leaf_55_clk),
    .D(net1938),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8410_ (.CLK(clknet_leaf_40_clk),
    .D(net1965),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8411_ (.CLK(clknet_leaf_61_clk),
    .D(net1924),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8412_ (.CLK(clknet_leaf_46_clk),
    .D(net1883),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8413_ (.CLK(clknet_leaf_61_clk),
    .D(net1896),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8414_ (.CLK(clknet_leaf_56_clk),
    .D(net1799),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8415_ (.CLK(clknet_leaf_51_clk),
    .D(net1906),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8416_ (.CLK(clknet_leaf_71_clk),
    .D(net1877),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8417_ (.CLK(clknet_leaf_69_clk),
    .D(net1813),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8418_ (.CLK(clknet_leaf_71_clk),
    .D(net1801),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8419_ (.CLK(clknet_leaf_55_clk),
    .D(net1889),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8420_ (.CLK(clknet_leaf_38_clk),
    .D(net981),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8421_ (.CLK(clknet_leaf_38_clk),
    .D(net1444),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8422_ (.CLK(clknet_leaf_38_clk),
    .D(net852),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8423_ (.CLK(clknet_leaf_32_clk),
    .D(net1572),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8424_ (.CLK(clknet_leaf_30_clk),
    .D(net1342),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8425_ (.CLK(clknet_leaf_19_clk),
    .D(net1159),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8426_ (.CLK(clknet_leaf_42_clk),
    .D(net1308),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8427_ (.CLK(clknet_leaf_68_clk),
    .D(net1015),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8428_ (.CLK(clknet_leaf_66_clk),
    .D(net1267),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8429_ (.CLK(clknet_leaf_41_clk),
    .D(net1352),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8430_ (.CLK(clknet_leaf_5_clk),
    .D(net1500),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8431_ (.CLK(clknet_leaf_71_clk),
    .D(net1422),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8432_ (.CLK(clknet_leaf_46_clk),
    .D(net1464),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8433_ (.CLK(clknet_leaf_41_clk),
    .D(net1279),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8434_ (.CLK(clknet_leaf_22_clk),
    .D(net1129),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8435_ (.CLK(clknet_leaf_26_clk),
    .D(net937),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8436_ (.CLK(clknet_leaf_51_clk),
    .D(net1606),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8437_ (.CLK(clknet_leaf_44_clk),
    .D(net1700),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8438_ (.CLK(clknet_leaf_20_clk),
    .D(net917),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8439_ (.CLK(clknet_leaf_29_clk),
    .D(net1512),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8440_ (.CLK(clknet_leaf_60_clk),
    .D(net959),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8441_ (.CLK(clknet_leaf_55_clk),
    .D(net1474),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8442_ (.CLK(clknet_leaf_40_clk),
    .D(net1470),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8443_ (.CLK(clknet_leaf_61_clk),
    .D(net1173),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8444_ (.CLK(clknet_leaf_31_clk),
    .D(net1586),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8445_ (.CLK(clknet_leaf_61_clk),
    .D(net1312),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8446_ (.CLK(clknet_leaf_56_clk),
    .D(net1428),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8447_ (.CLK(clknet_leaf_51_clk),
    .D(net1420),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8448_ (.CLK(clknet_leaf_71_clk),
    .D(net1759),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8449_ (.CLK(clknet_leaf_70_clk),
    .D(net1484),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8450_ (.CLK(clknet_leaf_70_clk),
    .D(net1466),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8451_ (.CLK(clknet_leaf_55_clk),
    .D(net1269),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8452_ (.CLK(clknet_leaf_36_clk),
    .D(net891),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8453_ (.CLK(clknet_leaf_32_clk),
    .D(net877),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8454_ (.CLK(clknet_leaf_36_clk),
    .D(net1053),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8455_ (.CLK(clknet_leaf_31_clk),
    .D(net879),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8456_ (.CLK(clknet_leaf_29_clk),
    .D(net1570),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8457_ (.CLK(clknet_leaf_19_clk),
    .D(net1201),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8458_ (.CLK(clknet_leaf_44_clk),
    .D(net1506),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8459_ (.CLK(clknet_leaf_71_clk),
    .D(net1235),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8460_ (.CLK(clknet_leaf_66_clk),
    .D(net1051),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8461_ (.CLK(clknet_leaf_45_clk),
    .D(net1482),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8462_ (.CLK(clknet_leaf_5_clk),
    .D(net1223),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8463_ (.CLK(clknet_leaf_71_clk),
    .D(net1318),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8464_ (.CLK(clknet_leaf_30_clk),
    .D(net1069),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8465_ (.CLK(clknet_leaf_45_clk),
    .D(net1324),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8466_ (.CLK(clknet_leaf_24_clk),
    .D(net1285),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8467_ (.CLK(clknet_leaf_10_clk),
    .D(net1518),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8468_ (.CLK(clknet_leaf_50_clk),
    .D(net1336),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8469_ (.CLK(clknet_leaf_47_clk),
    .D(net1123),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8470_ (.CLK(clknet_leaf_19_clk),
    .D(net1179),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8471_ (.CLK(clknet_leaf_32_clk),
    .D(net1003),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8472_ (.CLK(clknet_leaf_61_clk),
    .D(net1524),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8473_ (.CLK(clknet_leaf_57_clk),
    .D(net1450),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8474_ (.CLK(clknet_leaf_37_clk),
    .D(net1536),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8475_ (.CLK(clknet_leaf_62_clk),
    .D(net1702),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8476_ (.CLK(clknet_leaf_46_clk),
    .D(net1119),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8477_ (.CLK(clknet_leaf_69_clk),
    .D(net1300),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8478_ (.CLK(clknet_leaf_59_clk),
    .D(net1055),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8479_ (.CLK(clknet_leaf_50_clk),
    .D(net1291),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8480_ (.CLK(clknet_leaf_70_clk),
    .D(net1424),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8481_ (.CLK(clknet_leaf_69_clk),
    .D(net1382),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8482_ (.CLK(clknet_leaf_70_clk),
    .D(net1719),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8483_ (.CLK(clknet_leaf_58_clk),
    .D(net1789),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8484_ (.CLK(clknet_leaf_36_clk),
    .D(net1787),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8485_ (.CLK(clknet_leaf_36_clk),
    .D(net1775),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8486_ (.CLK(clknet_leaf_37_clk),
    .D(net1827),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8487_ (.CLK(clknet_leaf_31_clk),
    .D(net2130),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8488_ (.CLK(clknet_leaf_29_clk),
    .D(net1839),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8489_ (.CLK(clknet_leaf_25_clk),
    .D(net1898),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8490_ (.CLK(clknet_leaf_44_clk),
    .D(net1932),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8491_ (.CLK(clknet_leaf_69_clk),
    .D(net1887),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8492_ (.CLK(clknet_leaf_66_clk),
    .D(net1743),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8493_ (.CLK(clknet_leaf_41_clk),
    .D(net1912),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8494_ (.CLK(clknet_leaf_65_clk),
    .D(net1656),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8495_ (.CLK(clknet_leaf_67_clk),
    .D(net1618),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8496_ (.CLK(clknet_leaf_46_clk),
    .D(net1914),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8497_ (.CLK(clknet_leaf_41_clk),
    .D(net1908),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8498_ (.CLK(clknet_leaf_24_clk),
    .D(net1960),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8499_ (.CLK(clknet_leaf_26_clk),
    .D(net1660),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8500_ (.CLK(clknet_leaf_51_clk),
    .D(net1979),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8501_ (.CLK(clknet_leaf_44_clk),
    .D(net1962),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8502_ (.CLK(clknet_leaf_25_clk),
    .D(net1930),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8503_ (.CLK(clknet_leaf_32_clk),
    .D(net1944),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8504_ (.CLK(clknet_leaf_60_clk),
    .D(net1640),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8505_ (.CLK(clknet_leaf_56_clk),
    .D(net1771),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8506_ (.CLK(clknet_leaf_40_clk),
    .D(net1967),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8507_ (.CLK(clknet_leaf_61_clk),
    .D(net1845),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8508_ (.CLK(clknet_leaf_41_clk),
    .D(net1977),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8509_ (.CLK(clknet_leaf_61_clk),
    .D(net1869),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8510_ (.CLK(clknet_leaf_59_clk),
    .D(net1928),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8511_ (.CLK(clknet_leaf_51_clk),
    .D(net1981),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8512_ (.CLK(clknet_leaf_70_clk),
    .D(net1904),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8513_ (.CLK(clknet_leaf_69_clk),
    .D(net1809),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8514_ (.CLK(clknet_leaf_70_clk),
    .D(net1958),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8515_ (.CLK(clknet_leaf_54_clk),
    .D(net1863),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8516_ (.CLK(clknet_leaf_37_clk),
    .D(net911),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8517_ (.CLK(clknet_leaf_38_clk),
    .D(net865),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8518_ (.CLK(clknet_leaf_38_clk),
    .D(net889),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8519_ (.CLK(clknet_leaf_33_clk),
    .D(net1380),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8520_ (.CLK(clknet_leaf_32_clk),
    .D(net1213),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8521_ (.CLK(clknet_leaf_19_clk),
    .D(net1275),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8522_ (.CLK(clknet_leaf_43_clk),
    .D(net1163),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8523_ (.CLK(clknet_leaf_68_clk),
    .D(net1283),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8524_ (.CLK(clknet_leaf_5_clk),
    .D(net1468),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8525_ (.CLK(clknet_leaf_45_clk),
    .D(net1117),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8526_ (.CLK(clknet_leaf_5_clk),
    .D(net1584),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8527_ (.CLK(clknet_leaf_71_clk),
    .D(net1476),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8528_ (.CLK(clknet_leaf_30_clk),
    .D(net1101),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8529_ (.CLK(clknet_leaf_41_clk),
    .D(net1803),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8530_ (.CLK(clknet_leaf_20_clk),
    .D(net973),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8531_ (.CLK(clknet_leaf_16_clk),
    .D(net1522),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8532_ (.CLK(clknet_leaf_51_clk),
    .D(net1374),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8533_ (.CLK(clknet_leaf_47_clk),
    .D(net1346),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8534_ (.CLK(clknet_leaf_19_clk),
    .D(net1089),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8535_ (.CLK(clknet_leaf_27_clk),
    .D(net1356),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8536_ (.CLK(clknet_leaf_61_clk),
    .D(net1296),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8537_ (.CLK(clknet_leaf_57_clk),
    .D(net1384),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8538_ (.CLK(clknet_leaf_40_clk),
    .D(net1791),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8539_ (.CLK(clknet_leaf_61_clk),
    .D(net1418),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8540_ (.CLK(clknet_leaf_31_clk),
    .D(net1273),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8541_ (.CLK(clknet_leaf_69_clk),
    .D(net1127),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8542_ (.CLK(clknet_leaf_59_clk),
    .D(net1013),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8543_ (.CLK(clknet_leaf_51_clk),
    .D(net1731),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8544_ (.CLK(clknet_leaf_72_clk),
    .D(net999),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8545_ (.CLK(clknet_leaf_70_clk),
    .D(net1568),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8546_ (.CLK(clknet_leaf_73_clk),
    .D(net899),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8547_ (.CLK(clknet_leaf_54_clk),
    .D(net1322),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8548_ (.CLK(clknet_leaf_37_clk),
    .D(net1017),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8549_ (.CLK(clknet_leaf_35_clk),
    .D(net1011),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8550_ (.CLK(clknet_leaf_35_clk),
    .D(net951),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8551_ (.CLK(clknet_leaf_33_clk),
    .D(net1412),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8552_ (.CLK(clknet_leaf_32_clk),
    .D(net939),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8553_ (.CLK(clknet_leaf_19_clk),
    .D(net1408),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8554_ (.CLK(clknet_leaf_44_clk),
    .D(net1472),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8555_ (.CLK(clknet_leaf_68_clk),
    .D(net1147),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8556_ (.CLK(clknet_leaf_0_clk),
    .D(net1614),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8557_ (.CLK(clknet_leaf_45_clk),
    .D(net1193),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8558_ (.CLK(clknet_leaf_5_clk),
    .D(net1610),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8559_ (.CLK(clknet_leaf_72_clk),
    .D(net1113),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8560_ (.CLK(clknet_leaf_30_clk),
    .D(net1019),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8561_ (.CLK(clknet_leaf_41_clk),
    .D(net1662),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8562_ (.CLK(clknet_leaf_20_clk),
    .D(net955),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8563_ (.CLK(clknet_leaf_16_clk),
    .D(net1706),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8564_ (.CLK(clknet_leaf_51_clk),
    .D(net1544),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8565_ (.CLK(clknet_leaf_48_clk),
    .D(net1093),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8566_ (.CLK(clknet_leaf_19_clk),
    .D(net1364),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8567_ (.CLK(clknet_leaf_29_clk),
    .D(net1739),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8568_ (.CLK(clknet_leaf_61_clk),
    .D(net1372),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8569_ (.CLK(clknet_leaf_57_clk),
    .D(net1007),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8570_ (.CLK(clknet_leaf_40_clk),
    .D(net1446),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8571_ (.CLK(clknet_leaf_61_clk),
    .D(net1287),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8572_ (.CLK(clknet_leaf_31_clk),
    .D(net1227),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8573_ (.CLK(clknet_leaf_69_clk),
    .D(net1366),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8574_ (.CLK(clknet_leaf_59_clk),
    .D(net995),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8575_ (.CLK(clknet_leaf_51_clk),
    .D(net1582),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8576_ (.CLK(clknet_leaf_72_clk),
    .D(net1137),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8577_ (.CLK(clknet_leaf_70_clk),
    .D(net1765),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8578_ (.CLK(clknet_leaf_73_clk),
    .D(net967),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8579_ (.CLK(clknet_leaf_54_clk),
    .D(net1241),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ));
 sky130_fd_sc_hd__dfstp_1 _8580_ (.CLK(clknet_leaf_23_clk),
    .D(_1244_),
    .SET_B(_0260_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8581_ (.CLK(clknet_leaf_16_clk),
    .D(_1245_),
    .RESET_B(_0261_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8582_ (.CLK(clknet_leaf_16_clk),
    .D(_1246_),
    .RESET_B(_0262_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8583_ (.CLK(clknet_leaf_12_clk),
    .D(_1247_),
    .RESET_B(_0263_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8584_ (.CLK(clknet_leaf_11_clk),
    .D(_1248_),
    .RESET_B(_0264_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8585_ (.CLK(clknet_leaf_11_clk),
    .D(_1249_),
    .RESET_B(_0265_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8586_ (.CLK(clknet_leaf_13_clk),
    .D(_1250_),
    .RESET_B(_0266_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8587_ (.CLK(clknet_leaf_11_clk),
    .D(_1251_),
    .RESET_B(_0267_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8588_ (.CLK(clknet_leaf_3_clk),
    .D(_1252_),
    .RESET_B(_0268_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8589_ (.CLK(clknet_leaf_3_clk),
    .D(_1253_),
    .RESET_B(_0269_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8590_ (.CLK(clknet_leaf_13_clk),
    .D(_1254_),
    .RESET_B(_0270_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8591_ (.CLK(clknet_leaf_12_clk),
    .D(_1255_),
    .RESET_B(_0271_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8592_ (.CLK(clknet_leaf_15_clk),
    .D(net2029),
    .RESET_B(_0272_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8593_ (.CLK(clknet_leaf_15_clk),
    .D(net2018),
    .RESET_B(_0273_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8594_ (.CLK(clknet_leaf_10_clk),
    .D(_1258_),
    .RESET_B(_0274_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8595_ (.CLK(clknet_leaf_10_clk),
    .D(_1259_),
    .RESET_B(_0275_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8596_ (.CLK(clknet_leaf_22_clk),
    .D(net2032),
    .RESET_B(_0276_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8597_ (.CLK(clknet_leaf_22_clk),
    .D(_1261_),
    .RESET_B(_0277_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[19] ));
 sky130_fd_sc_hd__dfrtp_1 _8598_ (.CLK(clknet_leaf_22_clk),
    .D(_1262_),
    .RESET_B(_0278_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[20] ));
 sky130_fd_sc_hd__dfrtp_1 _8599_ (.CLK(clknet_leaf_49_clk),
    .D(_1263_),
    .RESET_B(_0279_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8600_ (.CLK(clknet_leaf_49_clk),
    .D(_1264_),
    .RESET_B(_0280_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8601_ (.CLK(clknet_leaf_49_clk),
    .D(_1265_),
    .RESET_B(_0281_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8602_ (.CLK(clknet_leaf_54_clk),
    .D(_1266_),
    .RESET_B(_0282_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8603_ (.CLK(clknet_leaf_58_clk),
    .D(_1267_),
    .RESET_B(_0283_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[25] ));
 sky130_fd_sc_hd__dfrtp_1 _8604_ (.CLK(clknet_leaf_58_clk),
    .D(_1268_),
    .RESET_B(_0284_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8605_ (.CLK(clknet_leaf_54_clk),
    .D(_1269_),
    .RESET_B(_0285_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[27] ));
 sky130_fd_sc_hd__dfrtp_1 _8606_ (.CLK(clknet_leaf_0_clk),
    .D(_1270_),
    .RESET_B(_0286_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[28] ));
 sky130_fd_sc_hd__dfrtp_1 _8607_ (.CLK(clknet_leaf_0_clk),
    .D(_1271_),
    .RESET_B(_0287_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[29] ));
 sky130_fd_sc_hd__dfrtp_1 _8608_ (.CLK(clknet_leaf_0_clk),
    .D(_1272_),
    .RESET_B(_0288_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[30] ));
 sky130_fd_sc_hd__dfrtp_1 _8609_ (.CLK(clknet_leaf_49_clk),
    .D(_1273_),
    .RESET_B(_0289_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8610_ (.CLK(clknet_leaf_37_clk),
    .D(net1761),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8611_ (.CLK(clknet_leaf_38_clk),
    .D(net2115),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8612_ (.CLK(clknet_leaf_35_clk),
    .D(net1879),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8613_ (.CLK(clknet_leaf_33_clk),
    .D(net1853),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8614_ (.CLK(clknet_leaf_29_clk),
    .D(net1934),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8615_ (.CLK(clknet_leaf_19_clk),
    .D(net2149),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8616_ (.CLK(clknet_leaf_44_clk),
    .D(net1849),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8617_ (.CLK(clknet_leaf_68_clk),
    .D(net1857),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8618_ (.CLK(clknet_leaf_5_clk),
    .D(net1971),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8619_ (.CLK(clknet_leaf_45_clk),
    .D(net1755),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8620_ (.CLK(clknet_leaf_4_clk),
    .D(net1841),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8621_ (.CLK(clknet_leaf_0_clk),
    .D(net1952),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8622_ (.CLK(clknet_leaf_30_clk),
    .D(net1668),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8623_ (.CLK(clknet_leaf_41_clk),
    .D(net1995),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8624_ (.CLK(clknet_leaf_25_clk),
    .D(net1910),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8625_ (.CLK(clknet_leaf_16_clk),
    .D(net1815),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8626_ (.CLK(clknet_leaf_50_clk),
    .D(net1936),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8627_ (.CLK(clknet_leaf_48_clk),
    .D(net1672),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8628_ (.CLK(clknet_leaf_20_clk),
    .D(net1715),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8629_ (.CLK(clknet_leaf_24_clk),
    .D(net1871),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8630_ (.CLK(clknet_leaf_61_clk),
    .D(net1821),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8631_ (.CLK(clknet_leaf_56_clk),
    .D(net1867),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8632_ (.CLK(clknet_leaf_40_clk),
    .D(net1833),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8633_ (.CLK(clknet_leaf_61_clk),
    .D(net1900),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8634_ (.CLK(clknet_leaf_31_clk),
    .D(net1807),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8635_ (.CLK(clknet_leaf_69_clk),
    .D(net1831),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8636_ (.CLK(clknet_leaf_60_clk),
    .D(net1598),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8637_ (.CLK(clknet_leaf_51_clk),
    .D(net1859),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8638_ (.CLK(clknet_leaf_72_clk),
    .D(net1634),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8639_ (.CLK(clknet_leaf_70_clk),
    .D(net1948),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8640_ (.CLK(clknet_leaf_73_clk),
    .D(net1410),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8641_ (.CLK(clknet_leaf_54_clk),
    .D(net1875),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8642_ (.CLK(clknet_leaf_40_clk),
    .D(net2047),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8643_ (.CLK(clknet_leaf_38_clk),
    .D(net1751),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8644_ (.CLK(clknet_leaf_38_clk),
    .D(net1793),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8645_ (.CLK(clknet_leaf_34_clk),
    .D(net1735),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8646_ (.CLK(clknet_leaf_29_clk),
    .D(net1785),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8647_ (.CLK(clknet_leaf_19_clk),
    .D(net2147),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8648_ (.CLK(clknet_leaf_43_clk),
    .D(net1835),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8649_ (.CLK(clknet_leaf_69_clk),
    .D(net1747),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8650_ (.CLK(clknet_leaf_5_clk),
    .D(net1946),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8651_ (.CLK(clknet_leaf_42_clk),
    .D(net1690),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8652_ (.CLK(clknet_leaf_4_clk),
    .D(net1767),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8653_ (.CLK(clknet_leaf_72_clk),
    .D(net1630),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8654_ (.CLK(clknet_leaf_46_clk),
    .D(net1783),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8655_ (.CLK(clknet_leaf_41_clk),
    .D(net1918),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8656_ (.CLK(clknet_leaf_25_clk),
    .D(net1861),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8657_ (.CLK(clknet_leaf_10_clk),
    .D(net1847),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8658_ (.CLK(clknet_leaf_52_clk),
    .D(net1855),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8659_ (.CLK(clknet_leaf_50_clk),
    .D(net1894),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8660_ (.CLK(clknet_leaf_21_clk),
    .D(net1779),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8661_ (.CLK(clknet_leaf_24_clk),
    .D(net1753),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8662_ (.CLK(clknet_leaf_60_clk),
    .D(net1763),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8663_ (.CLK(clknet_leaf_56_clk),
    .D(net1644),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8664_ (.CLK(clknet_leaf_40_clk),
    .D(net1865),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8665_ (.CLK(clknet_leaf_61_clk),
    .D(net1916),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8666_ (.CLK(clknet_leaf_31_clk),
    .D(net1817),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8667_ (.CLK(clknet_leaf_61_clk),
    .D(net1837),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8668_ (.CLK(clknet_leaf_56_clk),
    .D(net1749),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8669_ (.CLK(clknet_leaf_51_clk),
    .D(net1985),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8670_ (.CLK(clknet_leaf_72_clk),
    .D(net1708),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8671_ (.CLK(clknet_leaf_69_clk),
    .D(net1723),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8672_ (.CLK(clknet_leaf_70_clk),
    .D(net1922),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8673_ (.CLK(clknet_leaf_55_clk),
    .D(net1797),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8674_ (.CLK(clknet_leaf_6_clk),
    .D(_1338_),
    .Q(\U_DATAPATH.U_EX_MEM.i_result_src_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8675_ (.CLK(clknet_leaf_6_clk),
    .D(net2208),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8676_ (.CLK(clknet_leaf_6_clk),
    .D(_1340_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8677_ (.CLK(clknet_leaf_6_clk),
    .D(_1341_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8678_ (.CLK(clknet_leaf_6_clk),
    .D(_1342_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8679_ (.CLK(clknet_leaf_39_clk),
    .D(net921),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8680_ (.CLK(clknet_leaf_38_clk),
    .D(net1219),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8681_ (.CLK(clknet_leaf_38_clk),
    .D(net1496),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8682_ (.CLK(clknet_leaf_34_clk),
    .D(net1717),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8683_ (.CLK(clknet_leaf_30_clk),
    .D(net1378),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8684_ (.CLK(clknet_leaf_19_clk),
    .D(net1622),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8685_ (.CLK(clknet_leaf_43_clk),
    .D(net1073),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8686_ (.CLK(clknet_leaf_61_clk),
    .D(net1666),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8687_ (.CLK(clknet_leaf_5_clk),
    .D(net1628),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8688_ (.CLK(clknet_leaf_42_clk),
    .D(net1205),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8689_ (.CLK(clknet_leaf_6_clk),
    .D(net1546),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8690_ (.CLK(clknet_leaf_66_clk),
    .D(net1121),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8691_ (.CLK(clknet_leaf_46_clk),
    .D(net1534),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8692_ (.CLK(clknet_leaf_42_clk),
    .D(net1406),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8693_ (.CLK(clknet_leaf_25_clk),
    .D(net1652),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8694_ (.CLK(clknet_leaf_26_clk),
    .D(net1131),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8695_ (.CLK(clknet_leaf_52_clk),
    .D(net1632),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8696_ (.CLK(clknet_leaf_50_clk),
    .D(net1462),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8697_ (.CLK(clknet_leaf_21_clk),
    .D(net1081),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8698_ (.CLK(clknet_leaf_33_clk),
    .D(net1161),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8699_ (.CLK(clknet_leaf_60_clk),
    .D(net1530),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8700_ (.CLK(clknet_leaf_56_clk),
    .D(net1135),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8701_ (.CLK(clknet_leaf_40_clk),
    .D(net1532),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8702_ (.CLK(clknet_leaf_61_clk),
    .D(net1550),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8703_ (.CLK(clknet_leaf_37_clk),
    .D(net1578),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8704_ (.CLK(clknet_leaf_61_clk),
    .D(net1636),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8705_ (.CLK(clknet_leaf_57_clk),
    .D(net1257),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8706_ (.CLK(clknet_leaf_51_clk),
    .D(net1608),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8707_ (.CLK(clknet_leaf_71_clk),
    .D(net1488),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8708_ (.CLK(clknet_leaf_69_clk),
    .D(net1400),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8709_ (.CLK(clknet_leaf_70_clk),
    .D(net1670),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8710_ (.CLK(clknet_leaf_55_clk),
    .D(net1486),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8711_ (.CLK(clknet_leaf_65_clk),
    .D(_1375_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8712_ (.CLK(clknet_leaf_65_clk),
    .D(_1376_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8713_ (.CLK(clknet_leaf_65_clk),
    .D(_1377_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8714_ (.CLK(clknet_leaf_66_clk),
    .D(_1378_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8715_ (.CLK(clknet_leaf_48_clk),
    .D(_1379_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8716_ (.CLK(clknet_leaf_68_clk),
    .D(net2021),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8717_ (.CLK(clknet_leaf_62_clk),
    .D(net1294),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8718_ (.CLK(clknet_leaf_48_clk),
    .D(_1382_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8719_ (.CLK(clknet_leaf_63_clk),
    .D(_1383_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8720_ (.CLK(clknet_leaf_49_clk),
    .D(_1384_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8721_ (.CLK(clknet_leaf_63_clk),
    .D(_1385_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8722_ (.CLK(clknet_leaf_63_clk),
    .D(_1386_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8723_ (.CLK(clknet_leaf_29_clk),
    .D(net2107),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8724_ (.CLK(clknet_leaf_26_clk),
    .D(_1388_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8725_ (.CLK(clknet_leaf_28_clk),
    .D(net2183),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8726_ (.CLK(clknet_leaf_8_clk),
    .D(net2171),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8727_ (.CLK(clknet_leaf_9_clk),
    .D(net2145),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8728_ (.CLK(clknet_leaf_9_clk),
    .D(net2057),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8729_ (.CLK(clknet_leaf_9_clk),
    .D(net2094),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8730_ (.CLK(clknet_leaf_9_clk),
    .D(net2012),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8731_ (.CLK(clknet_leaf_9_clk),
    .D(_1395_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8732_ (.CLK(clknet_leaf_6_clk),
    .D(_1396_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8733_ (.CLK(clknet_leaf_6_clk),
    .D(_1397_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8734_ (.CLK(clknet_leaf_5_clk),
    .D(net2008),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8735_ (.CLK(clknet_leaf_6_clk),
    .D(_1399_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8736_ (.CLK(clknet_leaf_6_clk),
    .D(net1998),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8737_ (.CLK(clknet_leaf_6_clk),
    .D(_1401_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8738_ (.CLK(clknet_leaf_7_clk),
    .D(_1402_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8739_ (.CLK(clknet_leaf_25_clk),
    .D(_1403_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8740_ (.CLK(clknet_leaf_24_clk),
    .D(net2233),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8741_ (.CLK(clknet_leaf_27_clk),
    .D(_1405_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8742_ (.CLK(clknet_leaf_8_clk),
    .D(_1406_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[0] ));
 sky130_fd_sc_hd__ebufn_1 _8750_ (.A(net487),
    .TE_B(_3744_),
    .Z(_0064_));
 sky130_fd_sc_hd__conb_1 _8750__487 (.HI(net487));
 sky130_fd_sc_hd__ebufn_1 _8751_ (.A(net488),
    .TE_B(_3745_),
    .Z(_0065_));
 sky130_fd_sc_hd__conb_1 _8751__488 (.HI(net488));
 sky130_fd_sc_hd__ebufn_1 _8752_ (.A(net482),
    .TE_B(_3746_),
    .Z(_0066_));
 sky130_fd_sc_hd__conb_1 _8752__482 (.LO(net482));
 sky130_fd_sc_hd__ebufn_1 _8753_ (.A(net483),
    .TE_B(_3747_),
    .Z(_0067_));
 sky130_fd_sc_hd__conb_1 _8753__483 (.LO(net483));
 sky130_fd_sc_hd__ebufn_1 _8754_ (.A(net484),
    .TE_B(_3748_),
    .Z(_0068_));
 sky130_fd_sc_hd__conb_1 _8754__484 (.LO(net484));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__conb_1 core_485 (.LO(net485));
 sky130_fd_sc_hd__conb_1 core_486 (.LO(net486));
 sky130_fd_sc_hd__buf_6 fanout162 (.A(_2777_),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 fanout163 (.A(_2777_),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_8 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_8 fanout165 (.A(net170),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_8 fanout166 (.A(net170),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_8 fanout167 (.A(net169),
    .X(net167));
 sky130_fd_sc_hd__buf_8 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__buf_6 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_8 fanout170 (.A(_2652_),
    .X(net170));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(net174),
    .X(net171));
 sky130_fd_sc_hd__buf_4 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__buf_4 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 fanout174 (.A(_1910_),
    .X(net174));
 sky130_fd_sc_hd__buf_4 fanout175 (.A(net177),
    .X(net175));
 sky130_fd_sc_hd__buf_2 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__buf_4 fanout177 (.A(_1910_),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(net184),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 fanout180 (.A(net184),
    .X(net180));
 sky130_fd_sc_hd__buf_6 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__buf_6 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__buf_8 fanout184 (.A(_1910_),
    .X(net184));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 fanout186 (.A(_1721_),
    .X(net186));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_4 fanout188 (.A(_1721_),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_8 fanout189 (.A(net191),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__buf_4 fanout191 (.A(_1720_),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_8 fanout192 (.A(net194),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_8 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(_1698_),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_8 fanout195 (.A(_1698_),
    .X(net195));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(_1698_),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_8 fanout197 (.A(net199),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_8 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_8 fanout199 (.A(_1687_),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_8 fanout200 (.A(_1686_),
    .X(net200));
 sky130_fd_sc_hd__buf_4 fanout201 (.A(_1686_),
    .X(net201));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(_1672_),
    .X(net203));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(_1672_),
    .X(net204));
 sky130_fd_sc_hd__buf_4 fanout205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_8 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_4 fanout207 (.A(_1671_),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_8 fanout208 (.A(_1660_),
    .X(net208));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(_1660_),
    .X(net209));
 sky130_fd_sc_hd__buf_4 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 fanout211 (.A(_1660_),
    .X(net211));
 sky130_fd_sc_hd__buf_4 fanout212 (.A(_1659_),
    .X(net212));
 sky130_fd_sc_hd__buf_4 fanout213 (.A(_1659_),
    .X(net213));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(_1659_),
    .X(net214));
 sky130_fd_sc_hd__buf_8 fanout215 (.A(_3622_),
    .X(net215));
 sky130_fd_sc_hd__buf_8 fanout216 (.A(_3622_),
    .X(net216));
 sky130_fd_sc_hd__buf_8 fanout217 (.A(_3580_),
    .X(net217));
 sky130_fd_sc_hd__buf_6 fanout218 (.A(_3580_),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_16 fanout219 (.A(_3575_),
    .X(net219));
 sky130_fd_sc_hd__buf_6 fanout220 (.A(_3575_),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_8 fanout221 (.A(_2867_),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 fanout222 (.A(_2867_),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_8 fanout223 (.A(net225),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_8 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(_2866_),
    .X(net225));
 sky130_fd_sc_hd__buf_8 fanout226 (.A(_2774_),
    .X(net226));
 sky130_fd_sc_hd__buf_6 fanout227 (.A(_2774_),
    .X(net227));
 sky130_fd_sc_hd__buf_8 fanout228 (.A(_2770_),
    .X(net228));
 sky130_fd_sc_hd__buf_6 fanout229 (.A(_2770_),
    .X(net229));
 sky130_fd_sc_hd__buf_8 fanout230 (.A(_2765_),
    .X(net230));
 sky130_fd_sc_hd__buf_6 fanout231 (.A(_2765_),
    .X(net231));
 sky130_fd_sc_hd__buf_8 fanout232 (.A(_2761_),
    .X(net232));
 sky130_fd_sc_hd__buf_6 fanout233 (.A(_2761_),
    .X(net233));
 sky130_fd_sc_hd__buf_8 fanout234 (.A(_2756_),
    .X(net234));
 sky130_fd_sc_hd__buf_6 fanout235 (.A(_2756_),
    .X(net235));
 sky130_fd_sc_hd__buf_8 fanout236 (.A(_2750_),
    .X(net236));
 sky130_fd_sc_hd__buf_6 fanout237 (.A(_2750_),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_16 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__buf_12 fanout239 (.A(_3659_),
    .X(net239));
 sky130_fd_sc_hd__buf_8 fanout240 (.A(net241),
    .X(net240));
 sky130_fd_sc_hd__buf_12 fanout241 (.A(_3658_),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_16 fanout242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__buf_12 fanout243 (.A(_3625_),
    .X(net243));
 sky130_fd_sc_hd__buf_8 fanout244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_16 fanout245 (.A(_3624_),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_16 fanout246 (.A(_3620_),
    .X(net246));
 sky130_fd_sc_hd__buf_8 fanout247 (.A(_3620_),
    .X(net247));
 sky130_fd_sc_hd__buf_8 fanout248 (.A(_3618_),
    .X(net248));
 sky130_fd_sc_hd__buf_6 fanout249 (.A(_3618_),
    .X(net249));
 sky130_fd_sc_hd__buf_8 fanout250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__buf_12 fanout251 (.A(_3583_),
    .X(net251));
 sky130_fd_sc_hd__buf_8 fanout252 (.A(_3582_),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_8 fanout253 (.A(_3582_),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_16 fanout254 (.A(_3578_),
    .X(net254));
 sky130_fd_sc_hd__buf_6 fanout255 (.A(_3578_),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_16 fanout256 (.A(_3573_),
    .X(net256));
 sky130_fd_sc_hd__buf_8 fanout257 (.A(_3573_),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_16 fanout258 (.A(_3536_),
    .X(net258));
 sky130_fd_sc_hd__buf_8 fanout259 (.A(_3536_),
    .X(net259));
 sky130_fd_sc_hd__buf_8 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__buf_12 fanout261 (.A(_2772_),
    .X(net261));
 sky130_fd_sc_hd__buf_8 fanout262 (.A(_2768_),
    .X(net262));
 sky130_fd_sc_hd__buf_8 fanout263 (.A(_2768_),
    .X(net263));
 sky130_fd_sc_hd__buf_8 fanout264 (.A(_2763_),
    .X(net264));
 sky130_fd_sc_hd__buf_6 fanout265 (.A(_2763_),
    .X(net265));
 sky130_fd_sc_hd__buf_8 fanout266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_16 fanout267 (.A(_2759_),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_16 fanout268 (.A(_2754_),
    .X(net268));
 sky130_fd_sc_hd__buf_8 fanout269 (.A(_2754_),
    .X(net269));
 sky130_fd_sc_hd__buf_8 fanout270 (.A(_2748_),
    .X(net270));
 sky130_fd_sc_hd__buf_8 fanout271 (.A(_2748_),
    .X(net271));
 sky130_fd_sc_hd__buf_4 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__buf_4 fanout273 (.A(net281),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_4 fanout274 (.A(net281),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 fanout275 (.A(net281),
    .X(net275));
 sky130_fd_sc_hd__buf_4 fanout276 (.A(net281),
    .X(net276));
 sky130_fd_sc_hd__buf_4 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__buf_4 fanout279 (.A(net281),
    .X(net279));
 sky130_fd_sc_hd__buf_4 fanout280 (.A(net281),
    .X(net280));
 sky130_fd_sc_hd__buf_6 fanout281 (.A(_2206_),
    .X(net281));
 sky130_fd_sc_hd__buf_4 fanout282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__buf_2 fanout284 (.A(net292),
    .X(net284));
 sky130_fd_sc_hd__buf_4 fanout285 (.A(net292),
    .X(net285));
 sky130_fd_sc_hd__buf_2 fanout286 (.A(net292),
    .X(net286));
 sky130_fd_sc_hd__buf_4 fanout287 (.A(net292),
    .X(net287));
 sky130_fd_sc_hd__buf_4 fanout288 (.A(net290),
    .X(net288));
 sky130_fd_sc_hd__buf_4 fanout289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__buf_4 fanout290 (.A(net292),
    .X(net290));
 sky130_fd_sc_hd__buf_4 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__buf_4 fanout292 (.A(_2206_),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_8 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_8 fanout294 (.A(net298),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_8 fanout295 (.A(net298),
    .X(net295));
 sky130_fd_sc_hd__buf_4 fanout296 (.A(net297),
    .X(net296));
 sky130_fd_sc_hd__buf_4 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__buf_4 fanout298 (.A(_2205_),
    .X(net298));
 sky130_fd_sc_hd__buf_4 fanout299 (.A(_2205_),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_4 fanout300 (.A(_2205_),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_8 fanout301 (.A(net302),
    .X(net301));
 sky130_fd_sc_hd__buf_4 fanout302 (.A(_2205_),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_16 fanout304 (.A(_1466_),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_16 fanout305 (.A(_1466_),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_16 fanout306 (.A(_1464_),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_16 fanout307 (.A(_1464_),
    .X(net307));
 sky130_fd_sc_hd__buf_8 fanout308 (.A(_1447_),
    .X(net308));
 sky130_fd_sc_hd__buf_6 fanout309 (.A(_1447_),
    .X(net309));
 sky130_fd_sc_hd__buf_8 fanout310 (.A(_3616_),
    .X(net310));
 sky130_fd_sc_hd__buf_8 fanout311 (.A(_3616_),
    .X(net311));
 sky130_fd_sc_hd__buf_8 fanout312 (.A(net313),
    .X(net312));
 sky130_fd_sc_hd__buf_12 fanout313 (.A(_3540_),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_16 fanout314 (.A(_3539_),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_8 fanout315 (.A(_3539_),
    .X(net315));
 sky130_fd_sc_hd__buf_8 fanout316 (.A(net317),
    .X(net316));
 sky130_fd_sc_hd__buf_12 fanout317 (.A(_3534_),
    .X(net317));
 sky130_fd_sc_hd__buf_6 fanout319 (.A(_2861_),
    .X(net319));
 sky130_fd_sc_hd__buf_4 fanout320 (.A(_1834_),
    .X(net320));
 sky130_fd_sc_hd__buf_4 fanout321 (.A(_1821_),
    .X(net321));
 sky130_fd_sc_hd__buf_4 fanout322 (.A(_1810_),
    .X(net322));
 sky130_fd_sc_hd__buf_4 fanout323 (.A(_1800_),
    .X(net323));
 sky130_fd_sc_hd__buf_4 fanout324 (.A(_1788_),
    .X(net324));
 sky130_fd_sc_hd__buf_4 fanout325 (.A(_1777_),
    .X(net325));
 sky130_fd_sc_hd__buf_4 fanout326 (.A(_1767_),
    .X(net326));
 sky130_fd_sc_hd__buf_4 fanout327 (.A(_1757_),
    .X(net327));
 sky130_fd_sc_hd__buf_4 fanout328 (.A(_1728_),
    .X(net328));
 sky130_fd_sc_hd__buf_4 fanout329 (.A(_1716_),
    .X(net329));
 sky130_fd_sc_hd__buf_4 fanout330 (.A(_1707_),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_8 fanout331 (.A(_1695_),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_8 fanout332 (.A(_1679_),
    .X(net332));
 sky130_fd_sc_hd__buf_4 fanout333 (.A(_1667_),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_8 fanout334 (.A(_1655_),
    .X(net334));
 sky130_fd_sc_hd__buf_4 fanout335 (.A(_1643_),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_8 fanout336 (.A(_1630_),
    .X(net336));
 sky130_fd_sc_hd__buf_4 fanout337 (.A(_1619_),
    .X(net337));
 sky130_fd_sc_hd__buf_4 fanout338 (.A(_1607_),
    .X(net338));
 sky130_fd_sc_hd__buf_4 fanout339 (.A(_1595_),
    .X(net339));
 sky130_fd_sc_hd__buf_4 fanout340 (.A(_1584_),
    .X(net340));
 sky130_fd_sc_hd__buf_4 fanout341 (.A(_1572_),
    .X(net341));
 sky130_fd_sc_hd__buf_4 fanout342 (.A(_1562_),
    .X(net342));
 sky130_fd_sc_hd__buf_4 fanout343 (.A(_1550_),
    .X(net343));
 sky130_fd_sc_hd__buf_4 fanout344 (.A(_1537_),
    .X(net344));
 sky130_fd_sc_hd__buf_4 fanout345 (.A(_1526_),
    .X(net345));
 sky130_fd_sc_hd__buf_4 fanout346 (.A(_1496_),
    .X(net346));
 sky130_fd_sc_hd__buf_4 fanout347 (.A(_1485_),
    .X(net347));
 sky130_fd_sc_hd__buf_4 fanout348 (.A(_1473_),
    .X(net348));
 sky130_fd_sc_hd__buf_6 fanout349 (.A(_1457_),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_8 fanout350 (.A(_1457_),
    .X(net350));
 sky130_fd_sc_hd__buf_8 fanout351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_8 fanout353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_8 fanout354 (.A(_1431_),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_16 fanout355 (.A(_1430_),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_16 fanout356 (.A(net357),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_8 fanout358 (.A(_2863_),
    .X(net358));
 sky130_fd_sc_hd__buf_8 fanout359 (.A(net360),
    .X(net359));
 sky130_fd_sc_hd__buf_8 fanout360 (.A(_2860_),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_8 fanout361 (.A(net362),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_8 fanout362 (.A(_2857_),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_8 fanout363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_8 fanout364 (.A(_2856_),
    .X(net364));
 sky130_fd_sc_hd__buf_6 fanout366 (.A(_1453_),
    .X(net366));
 sky130_fd_sc_hd__buf_4 fanout367 (.A(_1453_),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_16 fanout368 (.A(_1471_),
    .X(net368));
 sky130_fd_sc_hd__buf_8 fanout369 (.A(_1471_),
    .X(net369));
 sky130_fd_sc_hd__buf_4 fanout370 (.A(_1446_),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_16 fanout371 (.A(_1445_),
    .X(net371));
 sky130_fd_sc_hd__buf_8 fanout372 (.A(_1445_),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_16 fanout373 (.A(_1444_),
    .X(net373));
 sky130_fd_sc_hd__buf_8 fanout374 (.A(_1444_),
    .X(net374));
 sky130_fd_sc_hd__buf_8 fanout375 (.A(_1414_),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_4 fanout376 (.A(_1414_),
    .X(net376));
 sky130_fd_sc_hd__buf_8 fanout377 (.A(net378),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_16 fanout378 (.A(\U_DATAPATH.U_ID_EX.o_addr_src_EX ),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_16 fanout379 (.A(net2315),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_8 fanout380 (.A(net2315),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_16 fanout381 (.A(net383),
    .X(net381));
 sky130_fd_sc_hd__buf_8 fanout382 (.A(net383),
    .X(net382));
 sky130_fd_sc_hd__buf_8 fanout383 (.A(net2167),
    .X(net383));
 sky130_fd_sc_hd__buf_8 fanout384 (.A(net385),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_16 fanout385 (.A(net2256),
    .X(net385));
 sky130_fd_sc_hd__buf_8 fanout386 (.A(net387),
    .X(net386));
 sky130_fd_sc_hd__buf_8 fanout387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_8 fanout388 (.A(net2256),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_8 fanout389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__buf_4 fanout390 (.A(net392),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_8 fanout391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__buf_8 fanout392 (.A(net398),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_8 fanout393 (.A(net398),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_8 fanout394 (.A(net397),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_8 fanout395 (.A(net396),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_8 fanout396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__buf_4 fanout397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__buf_8 fanout398 (.A(net2168),
    .X(net398));
 sky130_fd_sc_hd__buf_8 fanout399 (.A(net400),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_8 fanout400 (.A(net402),
    .X(net400));
 sky130_fd_sc_hd__buf_8 fanout401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_16 fanout402 (.A(net2166),
    .X(net402));
 sky130_fd_sc_hd__buf_8 fanout403 (.A(net408),
    .X(net403));
 sky130_fd_sc_hd__buf_8 fanout404 (.A(net407),
    .X(net404));
 sky130_fd_sc_hd__buf_8 fanout405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__buf_8 fanout406 (.A(net407),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_8 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_8 fanout408 (.A(net2166),
    .X(net408));
 sky130_fd_sc_hd__buf_8 fanout409 (.A(net2235),
    .X(net409));
 sky130_fd_sc_hd__buf_8 fanout410 (.A(net2235),
    .X(net410));
 sky130_fd_sc_hd__buf_6 fanout411 (.A(net413),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_4 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_8 fanout413 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ),
    .X(net413));
 sky130_fd_sc_hd__buf_6 fanout414 (.A(net416),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_8 fanout415 (.A(net416),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_8 fanout416 (.A(net2181),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_8 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_4 fanout418 (.A(net420),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_8 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__buf_8 fanout420 (.A(net426),
    .X(net420));
 sky130_fd_sc_hd__buf_6 fanout421 (.A(net426),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_8 fanout422 (.A(net425),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_8 fanout423 (.A(net424),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_8 fanout424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__buf_4 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__buf_8 fanout426 (.A(net2169),
    .X(net426));
 sky130_fd_sc_hd__buf_8 fanout427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_8 fanout428 (.A(net430),
    .X(net428));
 sky130_fd_sc_hd__buf_8 fanout429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_16 fanout430 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net430));
 sky130_fd_sc_hd__buf_8 fanout431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__buf_4 fanout432 (.A(net2143),
    .X(net432));
 sky130_fd_sc_hd__buf_8 fanout433 (.A(net436),
    .X(net433));
 sky130_fd_sc_hd__buf_8 fanout434 (.A(net436),
    .X(net434));
 sky130_fd_sc_hd__buf_4 fanout435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__buf_4 fanout436 (.A(net2143),
    .X(net436));
 sky130_fd_sc_hd__buf_8 fanout437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_16 fanout438 (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .X(net438));
 sky130_fd_sc_hd__buf_4 fanout439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_4 fanout440 (.A(net442),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_4 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_4 fanout442 (.A(net472),
    .X(net442));
 sky130_fd_sc_hd__buf_4 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__buf_4 fanout444 (.A(net472),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_4 fanout445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_4 fanout446 (.A(net472),
    .X(net446));
 sky130_fd_sc_hd__buf_4 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_4 fanout448 (.A(net454),
    .X(net448));
 sky130_fd_sc_hd__buf_4 fanout449 (.A(net454),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_4 fanout450 (.A(net454),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_2 fanout451 (.A(net454),
    .X(net451));
 sky130_fd_sc_hd__buf_4 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_4 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_8 fanout454 (.A(net472),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_4 fanout455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_4 fanout456 (.A(net459),
    .X(net456));
 sky130_fd_sc_hd__buf_4 fanout457 (.A(net459),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_4 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_4 fanout459 (.A(net472),
    .X(net459));
 sky130_fd_sc_hd__buf_4 fanout460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_4 fanout461 (.A(net472),
    .X(net461));
 sky130_fd_sc_hd__buf_4 fanout462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__buf_4 fanout463 (.A(net472),
    .X(net463));
 sky130_fd_sc_hd__buf_4 fanout464 (.A(net471),
    .X(net464));
 sky130_fd_sc_hd__buf_4 fanout465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_4 fanout466 (.A(net471),
    .X(net466));
 sky130_fd_sc_hd__buf_4 fanout467 (.A(net471),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_4 fanout468 (.A(net471),
    .X(net468));
 sky130_fd_sc_hd__buf_4 fanout469 (.A(net470),
    .X(net469));
 sky130_fd_sc_hd__buf_4 fanout470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_8 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__buf_8 fanout472 (.A(_0101_),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_16 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_8 fanout474 (.A(net475),
    .X(net474));
 sky130_fd_sc_hd__buf_6 fanout475 (.A(net63),
    .X(net475));
 sky130_fd_sc_hd__buf_6 fanout476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__buf_8 fanout477 (.A(net63),
    .X(net477));
 sky130_fd_sc_hd__buf_8 fanout478 (.A(net479),
    .X(net478));
 sky130_fd_sc_hd__buf_6 fanout479 (.A(net63),
    .X(net479));
 sky130_fd_sc_hd__buf_8 fanout480 (.A(net63),
    .X(net480));
 sky130_fd_sc_hd__buf_4 fanout481 (.A(net63),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[3] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[8] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(_1159_),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(_0506_),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(_1348_),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(_0423_),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(_0440_),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_0896_),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(_1351_),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(_1317_),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(_1359_),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(_1302_),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(_1368_),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[16] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(_1025_),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(_1168_),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(_0435_),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(_1327_),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(_0475_),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_0936_),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(_0596_),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(_0603_),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(_1357_),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(_0514_),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(_1158_),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[18] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(_0599_),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(_1163_),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(_1225_),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(_0494_),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(_1350_),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0938_),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(_1286_),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(_1373_),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(_1291_),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(_0446_),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(_1058_),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[4] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(_0578_),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(_0576_),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(_0601_),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(_0577_),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(_1072_),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0892_),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(_0560_),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(_1315_),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(_0600_),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(_0434_),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(_0412_),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[22] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(_0482_),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(_1101_),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(_1139_),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(_0588_),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(_1227_),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0942_),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(_1334_),
    .X(net1708));
 sky130_fd_sc_hd__buf_1 hold1092 (.A(net2110),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(_1064_),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(_0429_),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(_1292_),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0640_),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[18] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(_1346_),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(_1146_),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(_0573_),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(_1335_),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(_0418_),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0800_),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(_0500_),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(_1044_),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(_1207_),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(_0556_),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(_1309_),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[4] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(_0488_),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(_1231_),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(_0597_),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(_1156_),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(_0562_),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_0924_),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(_1313_),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(_1332_),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(_1307_),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(_1325_),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(_1283_),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\U_DATAPATH.U_EX_MEM.o_reg_write_M ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(_0493_),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(_1112_),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(_1274_),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(_1326_),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(_1241_),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0885_),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(_1316_),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(_1053_),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(_1169_),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(_1055_),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(_1149_),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[2] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(_1070_),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(_1324_),
    .X(net1779));
 sky130_fd_sc_hd__buf_1 hold1163 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[2] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(_0091_),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(_1318_),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(_1310_),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0784_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(_1148_),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(_1147_),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(_1202_),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(_1308_),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(_0589_),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[20] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(_1337_),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(_1078_),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(_1082_),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(_1193_),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(_0555_),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0340_),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(_1298_),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(_1177_),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[30] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(_0637_),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(_1081_),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(_1289_),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[14] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[5] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(_1330_),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(_0563_),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(_1294_),
    .X(net1821));
 sky130_fd_sc_hd__buf_1 hold1205 (.A(net2387),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(_0072_),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(_0595_),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_0893_),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(_1150_),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[21] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(_0341_),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(_1299_),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(_1296_),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(_1312_),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\U_DATAPATH.U_EX_MEM.i_funct3_EX[0] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(_1331_),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(_1152_),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(_1284_),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(_0540_),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(_1171_),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0882_),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(_1321_),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(_1280_),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[31] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(_0351_),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(_1277_),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(_1322_),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[2] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(_1281_),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(_1301_),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(_1320_),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(_1179_),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(_1328_),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_0890_),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(_1295_),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(_1173_),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(_1293_),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(_1052_),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(_1305_),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[24] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(_1080_),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(_1276_),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(_1063_),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(_1076_),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(_1069_),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_0806_),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(_1155_),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(_1083_),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(_1056_),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[18] ),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(_1323_),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(_1077_),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[7] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(_1153_),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(_1297_),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(_1057_),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(_1176_),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(_1079_),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0895_),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(_1161_),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(_1288_),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(_1157_),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(_1160_),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(_1329_),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0902_),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[12] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(_1319_),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[9] ),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(_0100_),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(_1336_),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(_1075_),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(_1067_),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_0794_),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(_1174_),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(_1166_),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(_1154_),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(_1278_),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(_1290_),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[9] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(_1073_),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(\U_DATAPATH.U_EX_MEM.i_reg_write_EX ),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(_0848_),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(_1071_),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(_1167_),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(_1314_),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_0791_),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(_1303_),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[12] ),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(_0332_),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(_1285_),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(_1061_),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(_1062_),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[3] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(_1178_),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(_1162_),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(_1165_),
    .X(net1962));
 sky130_fd_sc_hd__buf_1 hold1346 (.A(net2375),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(_1074_),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0891_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(_1170_),
    .X(net1967));
 sky130_fd_sc_hd__clkbuf_2 hold1351 (.A(net2109),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[7] ),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(_1282_),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(_1059_),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(_1060_),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[4] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(_1172_),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(_1164_),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(_1175_),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[6] ),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(_0326_),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(_1333_),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0786_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(_1068_),
    .X(net1987));
 sky130_fd_sc_hd__buf_1 hold1371 (.A(net2061),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(_1065_),
    .X(net1990));
 sky130_fd_sc_hd__buf_1 hold1374 (.A(net2385),
    .X(net1991));
 sky130_fd_sc_hd__buf_1 hold1375 (.A(net2374),
    .X(net1992));
 sky130_fd_sc_hd__buf_1 hold1376 (.A(net2383),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(_1287_),
    .X(net1995));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1379 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[11] ),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[16] ),
    .X(net755));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1380 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[26] ),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(_1400_),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(_0613_),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[9] ),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(_0329_),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[31] ),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(_1448_),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[5] ),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(_0325_),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_0798_),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_2 hold1390 (.A(net2384),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(_1398_),
    .X(net2008));
 sky130_fd_sc_hd__buf_1 hold1392 (.A(net2378),
    .X(net2009));
 sky130_fd_sc_hd__clkbuf_8 hold1393 (.A(net2206),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(_3734_),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(_1394_),
    .X(net2012));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1396 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[4] ),
    .X(net2013));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1397 (.A(_1943_),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(_2256_),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[22] ),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[15] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[11] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[15] ),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(_1257_),
    .X(net2018));
 sky130_fd_sc_hd__buf_2 hold1402 (.A(net2394),
    .X(net2019));
 sky130_fd_sc_hd__buf_4 hold1403 (.A(_3714_),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(_1380_),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[31] ),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(_2181_),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(_2182_),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[14] ),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(net126),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_0899_),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .X(net2027));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1411 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[14] ),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(_1256_),
    .X(net2029));
 sky130_fd_sc_hd__buf_1 hold1413 (.A(net2382),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(\U_DATAPATH.U_EX_MEM.i_result_src_EX[0] ),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(_1260_),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[8] ),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(_1980_),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[5] ),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(net129),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[5] ),
    .X(net759));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1420 (.A(net124),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[10] ),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(_0887_),
    .X(net2040));
 sky130_fd_sc_hd__buf_1 hold1424 (.A(net128),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[16] ),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[28] ),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[31] ),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[0] ),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(_1695_),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_0925_),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(_1306_),
    .X(net2047));
 sky130_fd_sc_hd__buf_1 hold1431 (.A(net2377),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[29] ),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[22] ),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(net108),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[3] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(net125),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[7] ),
    .X(net2054));
 sky130_fd_sc_hd__buf_4 hold1438 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(_3732_),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[10] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(_1392_),
    .X(net2057));
 sky130_fd_sc_hd__buf_2 hold1441 (.A(net2403),
    .X(net2058));
 sky130_fd_sc_hd__clkbuf_4 hold1442 (.A(_2265_),
    .X(net2059));
 sky130_fd_sc_hd__buf_1 hold1443 (.A(net2379),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[28] ),
    .X(net2109));
 sky130_fd_sc_hd__buf_1 hold1445 (.A(net2376),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(net127),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(net113),
    .X(net2064));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1448 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[23] ),
    .X(net2065));
 sky130_fd_sc_hd__buf_1 hold1449 (.A(net2389),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_0792_),
    .X(net762));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1450 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[17] ),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(net105),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(net106),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[30] ),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(net103),
    .X(net2071));
 sky130_fd_sc_hd__buf_1 hold1455 (.A(net2405),
    .X(net2072));
 sky130_fd_sc_hd__buf_1 hold1456 (.A(net2407),
    .X(net2073));
 sky130_fd_sc_hd__buf_4 hold1457 (.A(_2264_),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(net115),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(net118),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[22] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(net101),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(net122),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[17] ),
    .X(net2079));
 sky130_fd_sc_hd__clkbuf_4 hold1463 (.A(net110),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(net102),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(net121),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(net112),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[12] ),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(_1822_),
    .X(net2085));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1469 (.A(net2398),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0804_),
    .X(net764));
 sky130_fd_sc_hd__buf_1 hold1470 (.A(net2393),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(net114),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(net100),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(net111),
    .X(net2090));
 sky130_fd_sc_hd__buf_1 hold1474 (.A(net2386),
    .X(net2091));
 sky130_fd_sc_hd__clkbuf_8 hold1475 (.A(net2215),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(_3733_),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(_1393_),
    .X(net2094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(net117),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(net107),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[20] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(net119),
    .X(net2097));
 sky130_fd_sc_hd__buf_1 hold1481 (.A(net2392),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(net120),
    .X(net2099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(_0888_),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(net116),
    .X(net2102));
 sky130_fd_sc_hd__clkbuf_2 hold1486 (.A(net2397),
    .X(net2103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(net104),
    .X(net2104));
 sky130_fd_sc_hd__buf_2 hold1488 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[19] ),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(_3726_),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_0908_),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(_1387_),
    .X(net2107));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1491 (.A(\U_CONTROL_UNIT.i_jump_EX ),
    .X(net2108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[15] ),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[8] ),
    .X(net2373));
 sky130_fd_sc_hd__buf_4 hold1494 (.A(net180),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .X(net2112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(_0889_),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(_1275_),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(net109),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0935_),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[19] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(net123),
    .X(net2117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(_0886_),
    .X(net2119));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1503 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[3] ),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(_1657_),
    .X(net2121));
 sky130_fd_sc_hd__clkbuf_2 hold1505 (.A(net2381),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ),
    .X(net2123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(_2120_),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(_2132_),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(_2133_),
    .X(net2126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_0079_),
    .X(net768));
 sky130_fd_sc_hd__buf_1 hold1510 (.A(net2395),
    .X(net2127));
 sky130_fd_sc_hd__buf_2 hold1511 (.A(net2388),
    .X(net2128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ),
    .X(net2129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(_1151_),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[2] ),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(_0322_),
    .X(net2132));
 sky130_fd_sc_hd__buf_1 hold1516 (.A(net2396),
    .X(net2133));
 sky130_fd_sc_hd__clkbuf_2 hold1517 (.A(net2380),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[3] ),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[20] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(_1054_),
    .X(net2137));
 sky130_fd_sc_hd__clkbuf_4 hold1521 (.A(net2400),
    .X(net2138));
 sky130_fd_sc_hd__clkbuf_2 hold1522 (.A(net2373),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[20] ),
    .X(net2140));
 sky130_fd_sc_hd__buf_2 hold1524 (.A(_1586_),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[15] ),
    .X(net2142));
 sky130_fd_sc_hd__clkbuf_2 hold1526 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net2143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(_3731_),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(_1391_),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_0802_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(_1311_),
    .X(net2147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(_1279_),
    .X(net2149));
 sky130_fd_sc_hd__buf_1 hold1533 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[0] ),
    .X(net2150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(_1920_),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(_0749_),
    .X(net2152));
 sky130_fd_sc_hd__buf_1 hold1536 (.A(net2399),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(\U_CONTROL_UNIT.i_branch_EX ),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[17] ),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(_0866_),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[2] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[28] ),
    .X(net2157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(_1474_),
    .X(net2158));
 sky130_fd_sc_hd__buf_1 hold1542 (.A(net2391),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(_2083_),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(_2096_),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(_2097_),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[8] ),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(_1778_),
    .X(net2165));
 sky130_fd_sc_hd__clkbuf_4 hold1549 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_0922_),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ),
    .X(net2169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(_3730_),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(_1390_),
    .X(net2171));
 sky130_fd_sc_hd__buf_2 hold1555 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[24] ),
    .X(net2172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[10] ),
    .X(net2173));
 sky130_fd_sc_hd__clkbuf_2 hold1557 (.A(_1769_),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[6] ),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(_1730_),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[23] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(_1955_),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(_1968_),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(_1969_),
    .X(net2180));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1564 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(_3729_),
    .X(net2182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(_1389_),
    .X(net2183));
 sky130_fd_sc_hd__clkbuf_2 hold1567 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ),
    .X(net2184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(_1965_),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(_1977_),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_0805_),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(_1978_),
    .X(net2187));
 sky130_fd_sc_hd__clkbuf_2 hold1571 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(_1897_),
    .X(net2189));
 sky130_fd_sc_hd__buf_4 hold1573 (.A(net2404),
    .X(net2190));
 sky130_fd_sc_hd__buf_1 hold1574 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ),
    .X(net2191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(_1946_),
    .X(net2192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(_1958_),
    .X(net2193));
 sky130_fd_sc_hd__clkbuf_2 hold1577 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(_2791_),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[7] ),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[3] ),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_4 hold1580 (.A(net2402),
    .X(net2197));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1581 (.A(_2261_),
    .X(net2198));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1582 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[11] ),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(_2114_),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(_2115_),
    .X(net2202));
 sky130_fd_sc_hd__clkbuf_2 hold1586 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .X(net2203));
 sky130_fd_sc_hd__buf_1 hold1587 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[1] ),
    .X(net2204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[11] ),
    .X(net2205));
 sky130_fd_sc_hd__clkbuf_2 hold1589 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_0785_),
    .X(net776));
 sky130_fd_sc_hd__buf_1 hold1590 (.A(_3692_),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(_1339_),
    .X(net2208));
 sky130_fd_sc_hd__buf_1 hold1592 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ),
    .X(net2209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(_2055_),
    .X(net2210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(_2111_),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(_2123_),
    .X(net2213));
 sky130_fd_sc_hd__clkbuf_8 hold1597 (.A(net2406),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[28] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[26] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(_2129_),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(_2141_),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(_2142_),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[19] ),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[27] ),
    .X(net2221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(_1644_),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ),
    .X(net2223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(_2011_),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(_2022_),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(_2023_),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_0914_),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[28] ),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(_2156_),
    .X(net2228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(_2168_),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(_2169_),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[4] ),
    .X(net2231));
 sky130_fd_sc_hd__buf_1 hold1615 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .X(net2232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(_1404_),
    .X(net2233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .X(net2234));
 sky130_fd_sc_hd__buf_4 hold1618 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[29] ),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[15] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(_1497_),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ),
    .X(net2238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(_2093_),
    .X(net2239));
 sky130_fd_sc_hd__buf_2 hold1623 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .X(net2240));
 sky130_fd_sc_hd__buf_1 hold1624 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ),
    .X(net2241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(_2028_),
    .X(net2242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(_2041_),
    .X(net2243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(_2042_),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[9] ),
    .X(net2245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[25] ),
    .X(net2246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_0903_),
    .X(net780));
 sky130_fd_sc_hd__buf_1 hold1630 (.A(_1608_),
    .X(net2247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[18] ),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(_2065_),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(_2077_),
    .X(net2250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(_2078_),
    .X(net2251));
 sky130_fd_sc_hd__buf_1 hold1635 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ),
    .X(net2252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(_2047_),
    .X(net2253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(_2058_),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(_2059_),
    .X(net2255));
 sky130_fd_sc_hd__buf_2 hold1639 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ),
    .X(net2256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[13] ),
    .X(net781));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1640 (.A(\U_DATAPATH.U_ID_EX.o_addr_src_EX ),
    .X(net2257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(_2813_),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(_2173_),
    .X(net2260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(_2175_),
    .X(net2261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(_2176_),
    .X(net2262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(_1912_),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(_1914_),
    .X(net2265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(_1928_),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_0901_),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[23] ),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(_1596_),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ),
    .X(net2269));
 sky130_fd_sc_hd__buf_1 hold1653 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[10] ),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(_1993_),
    .X(net2271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[5] ),
    .X(net2272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1656 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(_1984_),
    .X(net2275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[26] ),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[6] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[19] ),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(_2072_),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ),
    .X(net2279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(_2038_),
    .X(net2280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[30] ),
    .X(net2281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(_2147_),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(_2159_),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[13] ),
    .X(net2285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ),
    .X(net2286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_0926_),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(_2019_),
    .X(net2287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(_2031_),
    .X(net2288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[11] ),
    .X(net2289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(_2000_),
    .X(net2290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(_2002_),
    .X(net2291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[14] ),
    .X(net2292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[18] ),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(_1937_),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[17] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ),
    .X(net2297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(_1499_),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(_1500_),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(_3501_),
    .X(net2300));
 sky130_fd_sc_hd__buf_1 hold1684 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ),
    .X(net2301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(_1974_),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[21] ),
    .X(net2303));
 sky130_fd_sc_hd__buf_1 hold1687 (.A(_1564_),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1688 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(_2138_),
    .X(net2306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_0905_),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[3] ),
    .X(net2307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(_1940_),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[23] ),
    .X(net2309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(_1601_),
    .X(net2310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(_3400_),
    .X(net2311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(_0837_),
    .X(net2312));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1696 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[16] ),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[22] ),
    .X(net2314));
 sky130_fd_sc_hd__clkbuf_2 hold1698 (.A(\U_DATAPATH.U_ID_EX.o_alu_src_EX ),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(_1591_),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0810_),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[19] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[2] ),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[28] ),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[8] ),
    .X(net2319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(_1783_),
    .X(net2320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[5] ),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(_0819_),
    .X(net2322));
 sky130_fd_sc_hd__buf_1 hold1706 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(_1520_),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(_0831_),
    .X(net2325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[0] ),
    .X(net2326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_0939_),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[25] ),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[27] ),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(_0841_),
    .X(net2329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[1] ),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ),
    .X(net2331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(_0820_),
    .X(net2332));
 sky130_fd_sc_hd__buf_1 hold1716 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ),
    .X(net2333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(_1675_),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(_0816_),
    .X(net2335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ),
    .X(net2336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\U_DATAPATH.U_EX_MEM.o_result_src_M[0] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1720 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[18] ),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(_0832_),
    .X(net2338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[10] ),
    .X(net2339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(_0824_),
    .X(net2340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[21] ),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(_0835_),
    .X(net2342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ),
    .X(net2343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1727 (.A(_1490_),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[15] ),
    .X(net2345));
 sky130_fd_sc_hd__clkbuf_2 hold1729 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_0290_),
    .X(net790));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1730 (.A(_2861_),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(_0823_),
    .X(net2348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1732 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ),
    .X(net2349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(_1828_),
    .X(net2350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ),
    .X(net2351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(_0840_),
    .X(net2352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[14] ),
    .X(net2353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1737 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .X(net2354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(_2870_),
    .X(net2355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(_0814_),
    .X(net2356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[31] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[7] ),
    .X(net2357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(_1712_),
    .X(net2358));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1742 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ),
    .X(net2359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(_2002_),
    .X(net2360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1744 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ),
    .X(net2361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1745 (.A(_1793_),
    .X(net2362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1746 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ),
    .X(net2363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1747 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ),
    .X(net2364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1748 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[3] ),
    .X(net2365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[19] ),
    .X(net2366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_0813_),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1750 (.A(_1531_),
    .X(net2367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(_0833_),
    .X(net2368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ),
    .X(net2369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1753 (.A(\U_DATAPATH.U_ID_EX.o_addr_src_EX ),
    .X(net2370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[4] ),
    .X(net2371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1755 (.A(_0818_),
    .X(net2372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1756 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[30] ),
    .X(net2374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[21] ),
    .X(net2375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[29] ),
    .X(net2376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1759 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[13] ),
    .X(net2377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[21] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1760 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[11] ),
    .X(net2378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1761 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[27] ),
    .X(net2379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1762 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[3] ),
    .X(net2380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1763 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[16] ),
    .X(net2381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1764 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[18] ),
    .X(net2382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1765 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[26] ),
    .X(net2383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1766 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[28] ),
    .X(net2384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1767 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[27] ),
    .X(net2385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1768 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[13] ),
    .X(net2386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1769 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[12] ),
    .X(net2387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_0803_),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1770 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[0] ),
    .X(net2388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1771 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[10] ),
    .X(net2389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1772 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[24] ),
    .X(net2390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1773 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[6] ),
    .X(net2391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1774 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[25] ),
    .X(net2392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1775 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[26] ),
    .X(net2393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1776 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[31] ),
    .X(net2394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1777 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[4] ),
    .X(net2395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1778 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[0] ),
    .X(net2396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1779 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[2] ),
    .X(net2397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[0] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1780 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[16] ),
    .X(net2398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1781 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[25] ),
    .X(net2399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1782 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[29] ),
    .X(net2400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1783 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[25] ),
    .X(net2401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1784 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ),
    .X(net2402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1785 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ),
    .X(net2403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1786 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ),
    .X(net2404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1787 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[24] ),
    .X(net2405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1788 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[27] ),
    .X(net2406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1789 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ),
    .X(net2407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_0920_),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[22] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[3] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_0923_),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[1] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_0921_),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[2] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_0609_),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[11] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_0793_),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[29] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_0917_),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0910_),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[25] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_0807_),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[19] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_0907_),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[17] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_0799_),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[21] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_0941_),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[25] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_0945_),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[12] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[5] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[29] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_0666_),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[14] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_0934_),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[19] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_0801_),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[29] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_0811_),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[6] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_0894_),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0787_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[9] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_0929_),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[25] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_0913_),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[17] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_0937_),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[13] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_0933_),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[10] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_0647_),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[26] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[29] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_0949_),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[27] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_0915_),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\U_DATAPATH.U_EX_MEM.i_mem_write_EX ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0881_),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[12] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_0649_),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[11] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_0648_),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_0946_),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[27] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_0947_),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\U_DATAPATH.U_EX_MEM.i_funct3_EX[2] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_0884_),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_1086_),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[6] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_0788_),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_0476_),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[8] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_1021_),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[19] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_0656_),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_0479_),
    .X(net862));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold246 (.A(net2390),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_1181_),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0790_),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_0541_),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[11] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_0618_),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[24] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_0631_),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_0543_),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[6] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_0643_),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[8] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_1117_),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_1119_),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[18] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_0655_),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[4] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_0641_),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[9] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_0646_),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[27] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0645_),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_0809_),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_1182_),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_1116_),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_0415_),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[5] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_0612_),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[8] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[28] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_0615_),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_1210_),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_0414_),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[10] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_0617_),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_0509_),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[20] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_0916_),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_0627_),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_0445_),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_1180_),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[23] ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_0660_),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_0542_),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_0900_),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[20] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_1102_),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_1026_),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_1343_),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[12] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_0619_),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_1020_),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[28] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_0940_),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_0665_),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[7] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_0644_),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_0545_),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[9] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_0616_),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_0487_),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[15] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_1099_),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_1216_),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_0520_),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[22] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_0629_),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[7] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_0614_),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[3] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_0797_),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_0610_),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_0484_),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_1214_),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_1038_),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_1226_),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[21] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[24] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_0658_),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_1104_),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[14] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_0621_),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[31] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_0668_),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[15] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_0622_),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_0944_),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_1242_),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_0433_),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_0511_),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(_1194_),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[13] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_0620_),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[20] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[24] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_0657_),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[5] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_0642_),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_1084_),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_0510_),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_0470_),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_0912_),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_0590_),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_0569_),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_0444_),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[4] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_0611_),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_1238_),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[28] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_0464_),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_1208_),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_0552_),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_1135_),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[25] ),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_0632_),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0948_),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_1233_),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_0529_),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(_1213_),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_1206_),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_1091_),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\U_DATAPATH.U_EX_MEM.i_funct3_EX[1] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[26] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_1212_),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_1224_),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[31] ),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_0638_),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_0574_),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_0465_),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[22] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0808_),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_0659_),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[29] ),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_0636_),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_0421_),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_0431_),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[14] ),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_0651_),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[10] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_0526_),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_1046_),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_0443_),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_0473_),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_1045_),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_0898_),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_0468_),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[24] ),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_0661_),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(_1124_),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_1118_),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_1142_),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[23] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_0593_),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_1048_),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_0547_),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_0419_),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_0533_),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0343_),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_1031_),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_1128_),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(_0428_),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(_1349_),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(_0452_),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[26] ),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[13] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_0633_),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(_0502_),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_1361_),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(_0534_),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(_0432_),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[23] ),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0795_),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_0630_),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(_1198_),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(_0483_),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(_1229_),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(_0564_),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[17] ),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[10] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(_0654_),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(_1040_),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(_1192_),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(_0441_),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(_0462_),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0930_),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_1023_),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[27] ),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_0634_),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_0463_),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(_1223_),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(_1027_),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_0883_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[14] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_1189_),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_1140_),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_1354_),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_1133_),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_0491_),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0796_),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_1205_),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(_1098_),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(_1358_),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[21] ),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_0628_),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_1364_),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[11] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_1240_),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_0447_),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[25] ),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_0662_),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_0424_),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_0517_),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0931_),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_1219_),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_0417_),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_0449_),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_1035_),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_0416_),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[24] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[28] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_1631_),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_1089_),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_1362_),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_1186_),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_1029_),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0635_),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_0549_),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_0459_),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[30] ),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_0667_),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_1107_),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_0557_),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_0497_),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_1134_),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_0572_),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_0550_),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_0466_),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_0783_),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_0438_),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_0499_),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_0523_),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_1221_),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_0413_),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[30] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_1030_),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0530_),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_1121_),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_0495_),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_1352_),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0950_),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_0548_),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[26] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_0663_),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[27] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(_0664_),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_1184_),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_0591_),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ),
    .X(net1216));
 sky130_fd_sc_hd__clkbuf_2 hold6 (.A(net2050),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[23] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_0457_),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_1344_),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_0460_),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(_1126_),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_0598_),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0943_),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_1236_),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_0544_),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_0566_),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_1042_),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_1123_),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[31] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_0513_),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_0539_),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_1243_),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_0554_),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_0454_),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0951_),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(_0448_),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(_0496_),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(_0536_),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(_0453_),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(_0518_),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_1369_),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(_0471_),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_0504_),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(_0455_),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(_0508_),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0781_),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_1092_),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(_1115_),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_0420_),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_1204_),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(_1185_),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[23] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_1041_),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(_1097_),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(_0477_),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_1187_),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(_1130_),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_0911_),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(_1235_),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(_0503_),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_1143_),
    .X(net1291));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold675 (.A(net2401),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(_3720_),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(_1381_),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(_1200_),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(_0565_),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(_1141_),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(_0469_),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(_0528_),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(_0507_),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0780_),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(_1090_),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(_0561_),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(_1109_),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(_0489_),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[19] ),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(_0626_),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_0093_),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[9] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(_1127_),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(_0559_),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(_1211_),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(_1129_),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(_0442_),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0897_),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(_1037_),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(_0480_),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[17] ),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(_0624_),
    .X(net1332));
 sky130_fd_sc_hd__clkbuf_2 hold716 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[19] ),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(_0339_),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(_1132_),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[13] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(_0558_),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(_1028_),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(_1088_),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(_1049_),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(_1197_),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0650_),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(_1039_),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(_0522_),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(_1093_),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(_0461_),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(_1199_),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[21] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[2] ),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(_0639_),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(_0546_),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(_0505_),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(_1230_),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(_1237_),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_0909_),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(_0580_),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(_0568_),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(_1232_),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(_1196_),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(_1034_),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[7] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(_1347_),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(_1183_),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(_1145_),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(_1201_),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(_1033_),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_0789_),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(_0583_),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(_0567_),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(_0584_),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(_0478_),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(_0602_),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[16] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(_0532_),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(_1372_),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(_0456_),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(_0472_),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(_1356_),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_0904_),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(_1217_),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(_1304_),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(_1215_),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(_0575_),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(_0501_),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[15] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[31] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(_1203_),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(_1111_),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(_1095_),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(_1144_),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(_1050_),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_0919_),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(_1110_),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(_0579_),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(_0474_),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(_0512_),
    .X(net1434));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold818 (.A(\U_DATAPATH.U_EX_MEM.i_result_src_EX[1] ),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(_0847_),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[30] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(_0586_),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(_0537_),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(_0498_),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(_1085_),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(_1234_),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_0812_),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(_0524_),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(_1137_),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(_0451_),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(_0570_),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(_0551_),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[16] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(_0426_),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(_1032_),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(_1360_),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(_1096_),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(_1114_),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_0653_),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(_1188_),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(_1106_),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(_1218_),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(_1105_),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(_1191_),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[12] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(_0527_),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(_0582_),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(_1125_),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(_1113_),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(_1374_),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_0932_),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(_1371_),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(_0553_),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(_0594_),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(_0587_),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(_1345_),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[7] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(_0516_),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(_1094_),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(_0492_),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(_0430_),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(_1122_),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0927_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[1] ),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(_1420_),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(_0436_),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(_1103_),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(_0485_),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(_1043_),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0652_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[30] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(_1131_),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(_0571_),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(_1195_),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(_1136_),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(_1024_),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_0918_),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(_0439_),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(_1363_),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(_1365_),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(_1355_),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(_1138_),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[8] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(_0531_),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(_1036_),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(_0458_),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(_1228_),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(_1353_),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0928_),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(_0581_),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(_1366_),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(_0467_),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(_0585_),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(_0525_),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[18] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(_1022_),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(_0422_),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(_0519_),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(_0515_),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(_0481_),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_0906_),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(_1209_),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(_1120_),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(_1087_),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(_0425_),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(_0490_),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[18] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(_1367_),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(_0535_),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(_1239_),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(_1190_),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(_1108_),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0625_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(_0592_),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(_1047_),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(_0521_),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(_1051_),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(_1066_),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\U_DATAPATH.U_EX_MEM.o_result_src_M[1] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(_1300_),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(_0427_),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(_0486_),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(_0437_),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(_1100_),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0291_),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(_1370_),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(_1222_),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(_0450_),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(_1220_),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(_0538_),
    .X(net1616));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(i_instr_ID[10]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(i_instr_ID[19]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(i_instr_ID[20]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(i_instr_ID[21]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(i_instr_ID[22]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(i_instr_ID[23]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(i_instr_ID[24]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(i_instr_ID[25]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(i_instr_ID[26]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(i_instr_ID[27]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(i_instr_ID[28]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(i_instr_ID[11]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(i_instr_ID[29]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(i_instr_ID[2]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(i_instr_ID[30]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(i_instr_ID[31]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(i_instr_ID[3]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(i_instr_ID[4]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(i_instr_ID[5]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(i_instr_ID[6]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(i_instr_ID[7]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(i_instr_ID[8]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(i_instr_ID[12]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(i_instr_ID[9]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(i_read_data_M[0]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(i_read_data_M[10]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(i_read_data_M[11]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(i_read_data_M[12]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(i_read_data_M[13]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(i_read_data_M[14]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(i_read_data_M[15]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(i_read_data_M[16]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(i_read_data_M[17]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(i_instr_ID[13]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input40 (.A(i_read_data_M[18]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(i_read_data_M[19]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(i_read_data_M[1]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(i_read_data_M[20]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(i_read_data_M[21]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(i_read_data_M[22]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(i_read_data_M[23]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(i_read_data_M[24]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(i_read_data_M[25]),
    .X(net48));
 sky130_fd_sc_hd__buf_4 input49 (.A(i_read_data_M[26]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input5 (.A(i_instr_ID[14]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input50 (.A(i_read_data_M[27]),
    .X(net50));
 sky130_fd_sc_hd__dlymetal6s2s_1 input51 (.A(i_read_data_M[28]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(i_read_data_M[29]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(i_read_data_M[2]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(i_read_data_M[30]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(i_read_data_M[31]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(i_read_data_M[3]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(i_read_data_M[4]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(i_read_data_M[5]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(i_read_data_M[6]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(i_instr_ID[15]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(i_read_data_M[7]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(i_read_data_M[8]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(i_read_data_M[9]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_8 input63 (.A(rst),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input7 (.A(i_instr_ID[16]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(i_instr_ID[17]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(i_instr_ID[18]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 max_cap303 (.A(_2205_),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_2 max_cap318 (.A(_3534_),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_4 max_cap352 (.A(_1440_),
    .X(net352));
 sky130_fd_sc_hd__buf_4 max_cap357 (.A(_1430_),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_2 max_cap365 (.A(_2744_),
    .X(net365));
 sky130_fd_sc_hd__buf_12 output100 (.A(net100),
    .X(o_pc_IF[10]));
 sky130_fd_sc_hd__buf_12 output101 (.A(net101),
    .X(o_pc_IF[11]));
 sky130_fd_sc_hd__buf_12 output102 (.A(net102),
    .X(o_pc_IF[12]));
 sky130_fd_sc_hd__buf_12 output103 (.A(net103),
    .X(o_pc_IF[13]));
 sky130_fd_sc_hd__buf_12 output104 (.A(net104),
    .X(o_pc_IF[14]));
 sky130_fd_sc_hd__buf_12 output105 (.A(net105),
    .X(o_pc_IF[15]));
 sky130_fd_sc_hd__buf_12 output106 (.A(net106),
    .X(o_pc_IF[16]));
 sky130_fd_sc_hd__buf_12 output107 (.A(net107),
    .X(o_pc_IF[17]));
 sky130_fd_sc_hd__buf_12 output108 (.A(net108),
    .X(o_pc_IF[18]));
 sky130_fd_sc_hd__buf_12 output109 (.A(net109),
    .X(o_pc_IF[19]));
 sky130_fd_sc_hd__buf_12 output110 (.A(net110),
    .X(o_pc_IF[20]));
 sky130_fd_sc_hd__buf_12 output111 (.A(net111),
    .X(o_pc_IF[21]));
 sky130_fd_sc_hd__buf_12 output112 (.A(net112),
    .X(o_pc_IF[22]));
 sky130_fd_sc_hd__buf_12 output113 (.A(net113),
    .X(o_pc_IF[23]));
 sky130_fd_sc_hd__buf_12 output114 (.A(net114),
    .X(o_pc_IF[24]));
 sky130_fd_sc_hd__buf_12 output115 (.A(net115),
    .X(o_pc_IF[25]));
 sky130_fd_sc_hd__buf_12 output116 (.A(net116),
    .X(o_pc_IF[26]));
 sky130_fd_sc_hd__buf_12 output117 (.A(net117),
    .X(o_pc_IF[27]));
 sky130_fd_sc_hd__buf_12 output118 (.A(net118),
    .X(o_pc_IF[28]));
 sky130_fd_sc_hd__buf_12 output119 (.A(net119),
    .X(o_pc_IF[29]));
 sky130_fd_sc_hd__buf_12 output120 (.A(net120),
    .X(o_pc_IF[2]));
 sky130_fd_sc_hd__buf_12 output121 (.A(net121),
    .X(o_pc_IF[30]));
 sky130_fd_sc_hd__buf_12 output122 (.A(net122),
    .X(o_pc_IF[31]));
 sky130_fd_sc_hd__buf_12 output123 (.A(net123),
    .X(o_pc_IF[3]));
 sky130_fd_sc_hd__buf_12 output124 (.A(net124),
    .X(o_pc_IF[4]));
 sky130_fd_sc_hd__buf_12 output125 (.A(net125),
    .X(o_pc_IF[5]));
 sky130_fd_sc_hd__buf_12 output126 (.A(net126),
    .X(o_pc_IF[6]));
 sky130_fd_sc_hd__buf_12 output127 (.A(net127),
    .X(o_pc_IF[7]));
 sky130_fd_sc_hd__buf_12 output128 (.A(net128),
    .X(o_pc_IF[8]));
 sky130_fd_sc_hd__buf_12 output129 (.A(net129),
    .X(o_pc_IF[9]));
 sky130_fd_sc_hd__buf_12 output130 (.A(net130),
    .X(o_write_data_M[0]));
 sky130_fd_sc_hd__buf_12 output131 (.A(net131),
    .X(o_write_data_M[10]));
 sky130_fd_sc_hd__buf_12 output132 (.A(net132),
    .X(o_write_data_M[11]));
 sky130_fd_sc_hd__buf_12 output133 (.A(net133),
    .X(o_write_data_M[12]));
 sky130_fd_sc_hd__buf_12 output134 (.A(net134),
    .X(o_write_data_M[13]));
 sky130_fd_sc_hd__buf_12 output135 (.A(net135),
    .X(o_write_data_M[14]));
 sky130_fd_sc_hd__buf_12 output136 (.A(net136),
    .X(o_write_data_M[15]));
 sky130_fd_sc_hd__buf_12 output137 (.A(net137),
    .X(o_write_data_M[16]));
 sky130_fd_sc_hd__buf_12 output138 (.A(net138),
    .X(o_write_data_M[17]));
 sky130_fd_sc_hd__buf_12 output139 (.A(net139),
    .X(o_write_data_M[18]));
 sky130_fd_sc_hd__buf_12 output140 (.A(net140),
    .X(o_write_data_M[19]));
 sky130_fd_sc_hd__buf_12 output141 (.A(net141),
    .X(o_write_data_M[1]));
 sky130_fd_sc_hd__buf_12 output142 (.A(net142),
    .X(o_write_data_M[20]));
 sky130_fd_sc_hd__buf_12 output143 (.A(net143),
    .X(o_write_data_M[21]));
 sky130_fd_sc_hd__buf_12 output144 (.A(net144),
    .X(o_write_data_M[22]));
 sky130_fd_sc_hd__buf_12 output145 (.A(net145),
    .X(o_write_data_M[23]));
 sky130_fd_sc_hd__buf_12 output146 (.A(net146),
    .X(o_write_data_M[24]));
 sky130_fd_sc_hd__buf_12 output147 (.A(net147),
    .X(o_write_data_M[25]));
 sky130_fd_sc_hd__buf_12 output148 (.A(net148),
    .X(o_write_data_M[26]));
 sky130_fd_sc_hd__buf_12 output149 (.A(net149),
    .X(o_write_data_M[27]));
 sky130_fd_sc_hd__buf_12 output150 (.A(net150),
    .X(o_write_data_M[28]));
 sky130_fd_sc_hd__buf_12 output151 (.A(net151),
    .X(o_write_data_M[29]));
 sky130_fd_sc_hd__buf_12 output152 (.A(net152),
    .X(o_write_data_M[2]));
 sky130_fd_sc_hd__buf_12 output153 (.A(net153),
    .X(o_write_data_M[30]));
 sky130_fd_sc_hd__buf_12 output154 (.A(net154),
    .X(o_write_data_M[31]));
 sky130_fd_sc_hd__buf_12 output155 (.A(net155),
    .X(o_write_data_M[3]));
 sky130_fd_sc_hd__buf_12 output156 (.A(net156),
    .X(o_write_data_M[4]));
 sky130_fd_sc_hd__buf_12 output157 (.A(net157),
    .X(o_write_data_M[5]));
 sky130_fd_sc_hd__buf_12 output158 (.A(net158),
    .X(o_write_data_M[6]));
 sky130_fd_sc_hd__buf_12 output159 (.A(net159),
    .X(o_write_data_M[7]));
 sky130_fd_sc_hd__buf_12 output160 (.A(net160),
    .X(o_write_data_M[8]));
 sky130_fd_sc_hd__buf_12 output161 (.A(net161),
    .X(o_write_data_M[9]));
 sky130_fd_sc_hd__buf_12 output64 (.A(net64),
    .X(o_data_addr_M[0]));
 sky130_fd_sc_hd__buf_12 output65 (.A(net65),
    .X(o_data_addr_M[10]));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(o_data_addr_M[11]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(o_data_addr_M[12]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(o_data_addr_M[13]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(o_data_addr_M[14]));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(o_data_addr_M[15]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(o_data_addr_M[16]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net72),
    .X(o_data_addr_M[17]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(o_data_addr_M[18]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(o_data_addr_M[19]));
 sky130_fd_sc_hd__buf_12 output75 (.A(net75),
    .X(o_data_addr_M[1]));
 sky130_fd_sc_hd__buf_12 output76 (.A(net76),
    .X(o_data_addr_M[20]));
 sky130_fd_sc_hd__buf_12 output77 (.A(net77),
    .X(o_data_addr_M[21]));
 sky130_fd_sc_hd__buf_12 output78 (.A(net78),
    .X(o_data_addr_M[22]));
 sky130_fd_sc_hd__buf_12 output79 (.A(net79),
    .X(o_data_addr_M[23]));
 sky130_fd_sc_hd__buf_12 output80 (.A(net80),
    .X(o_data_addr_M[24]));
 sky130_fd_sc_hd__buf_12 output81 (.A(net81),
    .X(o_data_addr_M[25]));
 sky130_fd_sc_hd__buf_12 output82 (.A(net82),
    .X(o_data_addr_M[26]));
 sky130_fd_sc_hd__buf_12 output83 (.A(net83),
    .X(o_data_addr_M[27]));
 sky130_fd_sc_hd__buf_12 output84 (.A(net84),
    .X(o_data_addr_M[28]));
 sky130_fd_sc_hd__buf_12 output85 (.A(net85),
    .X(o_data_addr_M[29]));
 sky130_fd_sc_hd__buf_12 output86 (.A(net86),
    .X(o_data_addr_M[2]));
 sky130_fd_sc_hd__buf_12 output87 (.A(net87),
    .X(o_data_addr_M[30]));
 sky130_fd_sc_hd__buf_12 output88 (.A(net88),
    .X(o_data_addr_M[31]));
 sky130_fd_sc_hd__buf_12 output89 (.A(net89),
    .X(o_data_addr_M[3]));
 sky130_fd_sc_hd__buf_12 output90 (.A(net90),
    .X(o_data_addr_M[4]));
 sky130_fd_sc_hd__buf_12 output91 (.A(net91),
    .X(o_data_addr_M[5]));
 sky130_fd_sc_hd__buf_12 output92 (.A(net92),
    .X(o_data_addr_M[6]));
 sky130_fd_sc_hd__buf_12 output93 (.A(net93),
    .X(o_data_addr_M[7]));
 sky130_fd_sc_hd__buf_12 output94 (.A(net94),
    .X(o_data_addr_M[8]));
 sky130_fd_sc_hd__buf_12 output95 (.A(net95),
    .X(o_data_addr_M[9]));
 sky130_fd_sc_hd__buf_12 output96 (.A(net96),
    .X(o_funct3_MEM[0]));
 sky130_fd_sc_hd__buf_12 output97 (.A(net97),
    .X(o_funct3_MEM[1]));
 sky130_fd_sc_hd__buf_12 output98 (.A(net98),
    .X(o_funct3_MEM[2]));
 sky130_fd_sc_hd__buf_12 output99 (.A(net99),
    .X(o_mem_write_M));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(_1539_),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_4 split1 (.A(net184),
    .X(net2044));
 assign o_pc_IF[0] = net485;
 assign o_pc_IF[1] = net486;
endmodule

