magic
tech sky130A
magscale 1 2
timestamp 1730775358
<< obsli1 >>
rect 2760 2703 77280 76721
<< obsm1 >>
rect 14 2388 79934 76968
<< metal2 >>
rect 662 78618 718 79418
rect 2594 78618 2650 79418
rect 4526 78618 4582 79418
rect 6458 78618 6514 79418
rect 8390 78618 8446 79418
rect 10322 78618 10378 79418
rect 12254 78618 12310 79418
rect 14186 78618 14242 79418
rect 16118 78618 16174 79418
rect 18050 78618 18106 79418
rect 19982 78618 20038 79418
rect 21914 78618 21970 79418
rect 23846 78618 23902 79418
rect 25778 78618 25834 79418
rect 27710 78618 27766 79418
rect 29642 78618 29698 79418
rect 31574 78618 31630 79418
rect 33506 78618 33562 79418
rect 35438 78618 35494 79418
rect 37370 78618 37426 79418
rect 39302 78618 39358 79418
rect 41234 78618 41290 79418
rect 43166 78618 43222 79418
rect 45098 78618 45154 79418
rect 47030 78618 47086 79418
rect 48962 78618 49018 79418
rect 50250 78618 50306 79418
rect 52182 78618 52238 79418
rect 54114 78618 54170 79418
rect 56046 78618 56102 79418
rect 57978 78618 58034 79418
rect 59910 78618 59966 79418
rect 61842 78618 61898 79418
rect 63774 78618 63830 79418
rect 65706 78618 65762 79418
rect 67638 78618 67694 79418
rect 69570 78618 69626 79418
rect 71502 78618 71558 79418
rect 73434 78618 73490 79418
rect 75366 78618 75422 79418
rect 77298 78618 77354 79418
rect 79230 78618 79286 79418
rect 18 0 74 800
rect 1306 0 1362 800
rect 3238 0 3294 800
rect 5170 0 5226 800
rect 7102 0 7158 800
rect 9034 0 9090 800
rect 10966 0 11022 800
rect 12898 0 12954 800
rect 14830 0 14886 800
rect 16762 0 16818 800
rect 18694 0 18750 800
rect 20626 0 20682 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 26422 0 26478 800
rect 28354 0 28410 800
rect 30286 0 30342 800
rect 32218 0 32274 800
rect 34150 0 34206 800
rect 36082 0 36138 800
rect 38014 0 38070 800
rect 39946 0 40002 800
rect 41878 0 41934 800
rect 43810 0 43866 800
rect 45742 0 45798 800
rect 47674 0 47730 800
rect 49606 0 49662 800
rect 51538 0 51594 800
rect 53470 0 53526 800
rect 55402 0 55458 800
rect 57334 0 57390 800
rect 59266 0 59322 800
rect 61198 0 61254 800
rect 62486 0 62542 800
rect 64418 0 64474 800
rect 66350 0 66406 800
rect 68282 0 68338 800
rect 70214 0 70270 800
rect 72146 0 72202 800
rect 74078 0 74134 800
rect 76010 0 76066 800
rect 77942 0 77998 800
rect 79874 0 79930 800
<< obsm2 >>
rect 20 78562 606 78690
rect 774 78562 2538 78690
rect 2706 78562 4470 78690
rect 4638 78562 6402 78690
rect 6570 78562 8334 78690
rect 8502 78562 10266 78690
rect 10434 78562 12198 78690
rect 12366 78562 14130 78690
rect 14298 78562 16062 78690
rect 16230 78562 17994 78690
rect 18162 78562 19926 78690
rect 20094 78562 21858 78690
rect 22026 78562 23790 78690
rect 23958 78562 25722 78690
rect 25890 78562 27654 78690
rect 27822 78562 29586 78690
rect 29754 78562 31518 78690
rect 31686 78562 33450 78690
rect 33618 78562 35382 78690
rect 35550 78562 37314 78690
rect 37482 78562 39246 78690
rect 39414 78562 41178 78690
rect 41346 78562 43110 78690
rect 43278 78562 45042 78690
rect 45210 78562 46974 78690
rect 47142 78562 48906 78690
rect 49074 78562 50194 78690
rect 50362 78562 52126 78690
rect 52294 78562 54058 78690
rect 54226 78562 55990 78690
rect 56158 78562 57922 78690
rect 58090 78562 59854 78690
rect 60022 78562 61786 78690
rect 61954 78562 63718 78690
rect 63886 78562 65650 78690
rect 65818 78562 67582 78690
rect 67750 78562 69514 78690
rect 69682 78562 71446 78690
rect 71614 78562 73378 78690
rect 73546 78562 75310 78690
rect 75478 78562 77242 78690
rect 77410 78562 79174 78690
rect 79342 78562 79928 78690
rect 20 856 79928 78562
rect 130 800 1250 856
rect 1418 800 3182 856
rect 3350 800 5114 856
rect 5282 800 7046 856
rect 7214 800 8978 856
rect 9146 800 10910 856
rect 11078 800 12842 856
rect 13010 800 14774 856
rect 14942 800 16706 856
rect 16874 800 18638 856
rect 18806 800 20570 856
rect 20738 800 22502 856
rect 22670 800 24434 856
rect 24602 800 26366 856
rect 26534 800 28298 856
rect 28466 800 30230 856
rect 30398 800 32162 856
rect 32330 800 34094 856
rect 34262 800 36026 856
rect 36194 800 37958 856
rect 38126 800 39890 856
rect 40058 800 41822 856
rect 41990 800 43754 856
rect 43922 800 45686 856
rect 45854 800 47618 856
rect 47786 800 49550 856
rect 49718 800 51482 856
rect 51650 800 53414 856
rect 53582 800 55346 856
rect 55514 800 57278 856
rect 57446 800 59210 856
rect 59378 800 61142 856
rect 61310 800 62430 856
rect 62598 800 64362 856
rect 64530 800 66294 856
rect 66462 800 68226 856
rect 68394 800 70158 856
rect 70326 800 72090 856
rect 72258 800 74022 856
rect 74190 800 75954 856
rect 76122 800 77886 856
rect 78054 800 79818 856
<< metal3 >>
rect 0 78208 800 78328
rect 79242 78208 80042 78328
rect 0 76168 800 76288
rect 79242 76168 80042 76288
rect 0 74128 800 74248
rect 79242 74128 80042 74248
rect 0 72088 800 72208
rect 79242 72088 80042 72208
rect 0 70048 800 70168
rect 79242 70048 80042 70168
rect 0 68008 800 68128
rect 79242 68008 80042 68128
rect 0 65968 800 66088
rect 79242 65968 80042 66088
rect 0 64608 800 64728
rect 79242 63928 80042 64048
rect 0 62568 800 62688
rect 79242 61888 80042 62008
rect 0 60528 800 60648
rect 79242 59848 80042 59968
rect 0 58488 800 58608
rect 79242 57808 80042 57928
rect 0 56448 800 56568
rect 79242 55768 80042 55888
rect 0 54408 800 54528
rect 79242 53728 80042 53848
rect 0 52368 800 52488
rect 79242 51688 80042 51808
rect 0 50328 800 50448
rect 79242 49648 80042 49768
rect 0 48288 800 48408
rect 79242 47608 80042 47728
rect 0 46248 800 46368
rect 79242 46248 80042 46368
rect 0 44208 800 44328
rect 79242 44208 80042 44328
rect 0 42168 800 42288
rect 79242 42168 80042 42288
rect 0 40128 800 40248
rect 79242 40128 80042 40248
rect 0 38088 800 38208
rect 79242 38088 80042 38208
rect 0 36048 800 36168
rect 79242 36048 80042 36168
rect 0 34008 800 34128
rect 79242 34008 80042 34128
rect 0 31968 800 32088
rect 79242 31968 80042 32088
rect 0 29928 800 30048
rect 79242 29928 80042 30048
rect 0 27888 800 28008
rect 79242 27888 80042 28008
rect 0 25848 800 25968
rect 79242 25848 80042 25968
rect 0 23808 800 23928
rect 79242 23808 80042 23928
rect 0 21768 800 21888
rect 79242 21768 80042 21888
rect 0 19728 800 19848
rect 79242 19728 80042 19848
rect 0 17688 800 17808
rect 79242 17688 80042 17808
rect 0 15648 800 15768
rect 79242 15648 80042 15768
rect 0 13608 800 13728
rect 79242 13608 80042 13728
rect 0 11568 800 11688
rect 79242 11568 80042 11688
rect 0 9528 800 9648
rect 79242 9528 80042 9648
rect 0 7488 800 7608
rect 79242 7488 80042 7608
rect 0 5448 800 5568
rect 79242 5448 80042 5568
rect 0 3408 800 3528
rect 79242 3408 80042 3528
rect 0 1368 800 1488
rect 79242 1368 80042 1488
<< obsm3 >>
rect 880 78128 79162 78301
rect 800 76368 79242 78128
rect 880 76088 79162 76368
rect 800 74328 79242 76088
rect 880 74048 79162 74328
rect 800 72288 79242 74048
rect 880 72008 79162 72288
rect 800 70248 79242 72008
rect 880 69968 79162 70248
rect 800 68208 79242 69968
rect 880 67928 79162 68208
rect 800 66168 79242 67928
rect 880 65888 79162 66168
rect 800 64808 79242 65888
rect 880 64528 79242 64808
rect 800 64128 79242 64528
rect 800 63848 79162 64128
rect 800 62768 79242 63848
rect 880 62488 79242 62768
rect 800 62088 79242 62488
rect 800 61808 79162 62088
rect 800 60728 79242 61808
rect 880 60448 79242 60728
rect 800 60048 79242 60448
rect 800 59768 79162 60048
rect 800 58688 79242 59768
rect 880 58408 79242 58688
rect 800 58008 79242 58408
rect 800 57728 79162 58008
rect 800 56648 79242 57728
rect 880 56368 79242 56648
rect 800 55968 79242 56368
rect 800 55688 79162 55968
rect 800 54608 79242 55688
rect 880 54328 79242 54608
rect 800 53928 79242 54328
rect 800 53648 79162 53928
rect 800 52568 79242 53648
rect 880 52288 79242 52568
rect 800 51888 79242 52288
rect 800 51608 79162 51888
rect 800 50528 79242 51608
rect 880 50248 79242 50528
rect 800 49848 79242 50248
rect 800 49568 79162 49848
rect 800 48488 79242 49568
rect 880 48208 79242 48488
rect 800 47808 79242 48208
rect 800 47528 79162 47808
rect 800 46448 79242 47528
rect 880 46168 79162 46448
rect 800 44408 79242 46168
rect 880 44128 79162 44408
rect 800 42368 79242 44128
rect 880 42088 79162 42368
rect 800 40328 79242 42088
rect 880 40048 79162 40328
rect 800 38288 79242 40048
rect 880 38008 79162 38288
rect 800 36248 79242 38008
rect 880 35968 79162 36248
rect 800 34208 79242 35968
rect 880 33928 79162 34208
rect 800 32168 79242 33928
rect 880 31888 79162 32168
rect 800 30128 79242 31888
rect 880 29848 79162 30128
rect 800 28088 79242 29848
rect 880 27808 79162 28088
rect 800 26048 79242 27808
rect 880 25768 79162 26048
rect 800 24008 79242 25768
rect 880 23728 79162 24008
rect 800 21968 79242 23728
rect 880 21688 79162 21968
rect 800 19928 79242 21688
rect 880 19648 79162 19928
rect 800 17888 79242 19648
rect 880 17608 79162 17888
rect 800 15848 79242 17608
rect 880 15568 79162 15848
rect 800 13808 79242 15568
rect 880 13528 79162 13808
rect 800 11768 79242 13528
rect 880 11488 79162 11768
rect 800 9728 79242 11488
rect 880 9448 79162 9728
rect 800 7688 79242 9448
rect 880 7408 79162 7688
rect 800 5648 79242 7408
rect 880 5368 79162 5648
rect 800 3608 79242 5368
rect 880 3328 79162 3608
rect 800 1568 79242 3328
rect 880 1395 79162 1568
<< metal4 >>
rect 5864 2672 6184 76752
rect 6524 2672 6844 76752
rect 36584 2672 36904 76752
rect 37244 2672 37564 76752
rect 67304 2672 67624 76752
rect 67964 2672 68284 76752
<< obsm4 >>
rect 3187 3027 5784 76533
rect 6264 3027 6444 76533
rect 6924 3027 36504 76533
rect 36984 3027 37164 76533
rect 37644 3027 67224 76533
rect 67704 3027 67884 76533
rect 68364 3027 75565 76533
<< labels >>
rlabel metal2 s 62486 0 62542 800 6 clk
port 1 nsew signal input
rlabel metal2 s 39302 78618 39358 79418 6 i_instr_ID[0]
port 2 nsew signal input
rlabel metal3 s 79242 76168 80042 76288 6 i_instr_ID[10]
port 3 nsew signal input
rlabel metal3 s 79242 63928 80042 64048 6 i_instr_ID[11]
port 4 nsew signal input
rlabel metal2 s 47030 78618 47086 79418 6 i_instr_ID[12]
port 5 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 i_instr_ID[13]
port 6 nsew signal input
rlabel metal2 s 71502 78618 71558 79418 6 i_instr_ID[14]
port 7 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 i_instr_ID[15]
port 8 nsew signal input
rlabel metal3 s 79242 1368 80042 1488 6 i_instr_ID[16]
port 9 nsew signal input
rlabel metal2 s 48962 78618 49018 79418 6 i_instr_ID[17]
port 10 nsew signal input
rlabel metal3 s 79242 21768 80042 21888 6 i_instr_ID[18]
port 11 nsew signal input
rlabel metal3 s 79242 44208 80042 44328 6 i_instr_ID[19]
port 12 nsew signal input
rlabel metal2 s 27710 78618 27766 79418 6 i_instr_ID[1]
port 13 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 i_instr_ID[20]
port 14 nsew signal input
rlabel metal2 s 35438 78618 35494 79418 6 i_instr_ID[21]
port 15 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 i_instr_ID[22]
port 16 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 i_instr_ID[23]
port 17 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 i_instr_ID[24]
port 18 nsew signal input
rlabel metal3 s 79242 36048 80042 36168 6 i_instr_ID[25]
port 19 nsew signal input
rlabel metal2 s 8390 78618 8446 79418 6 i_instr_ID[26]
port 20 nsew signal input
rlabel metal2 s 54114 78618 54170 79418 6 i_instr_ID[27]
port 21 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 i_instr_ID[28]
port 22 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 i_instr_ID[29]
port 23 nsew signal input
rlabel metal2 s 79230 78618 79286 79418 6 i_instr_ID[2]
port 24 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 i_instr_ID[30]
port 25 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 i_instr_ID[31]
port 26 nsew signal input
rlabel metal3 s 79242 7488 80042 7608 6 i_instr_ID[3]
port 27 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 i_instr_ID[4]
port 28 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 i_instr_ID[5]
port 29 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 i_instr_ID[6]
port 30 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 i_instr_ID[7]
port 31 nsew signal input
rlabel metal2 s 21914 78618 21970 79418 6 i_instr_ID[8]
port 32 nsew signal input
rlabel metal2 s 45098 78618 45154 79418 6 i_instr_ID[9]
port 33 nsew signal input
rlabel metal2 s 73434 78618 73490 79418 6 i_read_data_M[0]
port 34 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 i_read_data_M[10]
port 35 nsew signal input
rlabel metal2 s 10322 78618 10378 79418 6 i_read_data_M[11]
port 36 nsew signal input
rlabel metal3 s 79242 61888 80042 62008 6 i_read_data_M[12]
port 37 nsew signal input
rlabel metal2 s 77298 78618 77354 79418 6 i_read_data_M[13]
port 38 nsew signal input
rlabel metal3 s 79242 57808 80042 57928 6 i_read_data_M[14]
port 39 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 i_read_data_M[15]
port 40 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 i_read_data_M[16]
port 41 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 i_read_data_M[17]
port 42 nsew signal input
rlabel metal3 s 79242 31968 80042 32088 6 i_read_data_M[18]
port 43 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 i_read_data_M[19]
port 44 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 i_read_data_M[1]
port 45 nsew signal input
rlabel metal3 s 79242 3408 80042 3528 6 i_read_data_M[20]
port 46 nsew signal input
rlabel metal2 s 31574 78618 31630 79418 6 i_read_data_M[21]
port 47 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 i_read_data_M[22]
port 48 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 i_read_data_M[23]
port 49 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 i_read_data_M[24]
port 50 nsew signal input
rlabel metal2 s 37370 78618 37426 79418 6 i_read_data_M[25]
port 51 nsew signal input
rlabel metal2 s 6458 78618 6514 79418 6 i_read_data_M[26]
port 52 nsew signal input
rlabel metal3 s 79242 59848 80042 59968 6 i_read_data_M[27]
port 53 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 i_read_data_M[28]
port 54 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 i_read_data_M[29]
port 55 nsew signal input
rlabel metal2 s 29642 78618 29698 79418 6 i_read_data_M[2]
port 56 nsew signal input
rlabel metal3 s 79242 17688 80042 17808 6 i_read_data_M[30]
port 57 nsew signal input
rlabel metal3 s 79242 68008 80042 68128 6 i_read_data_M[31]
port 58 nsew signal input
rlabel metal3 s 79242 25848 80042 25968 6 i_read_data_M[3]
port 59 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 i_read_data_M[4]
port 60 nsew signal input
rlabel metal3 s 79242 9528 80042 9648 6 i_read_data_M[5]
port 61 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 i_read_data_M[6]
port 62 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 i_read_data_M[7]
port 63 nsew signal input
rlabel metal3 s 79242 72088 80042 72208 6 i_read_data_M[8]
port 64 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 i_read_data_M[9]
port 65 nsew signal input
rlabel metal2 s 75366 78618 75422 79418 6 o_data_addr_M[0]
port 66 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 o_data_addr_M[10]
port 67 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 o_data_addr_M[11]
port 68 nsew signal output
rlabel metal2 s 56046 78618 56102 79418 6 o_data_addr_M[12]
port 69 nsew signal output
rlabel metal2 s 52182 78618 52238 79418 6 o_data_addr_M[13]
port 70 nsew signal output
rlabel metal2 s 25778 78618 25834 79418 6 o_data_addr_M[14]
port 71 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 o_data_addr_M[15]
port 72 nsew signal output
rlabel metal2 s 4526 78618 4582 79418 6 o_data_addr_M[16]
port 73 nsew signal output
rlabel metal3 s 79242 70048 80042 70168 6 o_data_addr_M[17]
port 74 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 o_data_addr_M[18]
port 75 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 o_data_addr_M[19]
port 76 nsew signal output
rlabel metal3 s 79242 55768 80042 55888 6 o_data_addr_M[1]
port 77 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 o_data_addr_M[20]
port 78 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 o_data_addr_M[21]
port 79 nsew signal output
rlabel metal3 s 79242 47608 80042 47728 6 o_data_addr_M[22]
port 80 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 o_data_addr_M[23]
port 81 nsew signal output
rlabel metal3 s 79242 15648 80042 15768 6 o_data_addr_M[24]
port 82 nsew signal output
rlabel metal2 s 19982 78618 20038 79418 6 o_data_addr_M[25]
port 83 nsew signal output
rlabel metal3 s 79242 29928 80042 30048 6 o_data_addr_M[26]
port 84 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 o_data_addr_M[27]
port 85 nsew signal output
rlabel metal2 s 69570 78618 69626 79418 6 o_data_addr_M[28]
port 86 nsew signal output
rlabel metal3 s 79242 34008 80042 34128 6 o_data_addr_M[29]
port 87 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 o_data_addr_M[2]
port 88 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 o_data_addr_M[30]
port 89 nsew signal output
rlabel metal2 s 50250 78618 50306 79418 6 o_data_addr_M[31]
port 90 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 o_data_addr_M[3]
port 91 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 o_data_addr_M[4]
port 92 nsew signal output
rlabel metal2 s 2594 78618 2650 79418 6 o_data_addr_M[5]
port 93 nsew signal output
rlabel metal2 s 12254 78618 12310 79418 6 o_data_addr_M[6]
port 94 nsew signal output
rlabel metal2 s 61842 78618 61898 79418 6 o_data_addr_M[7]
port 95 nsew signal output
rlabel metal2 s 63774 78618 63830 79418 6 o_data_addr_M[8]
port 96 nsew signal output
rlabel metal2 s 59910 78618 59966 79418 6 o_data_addr_M[9]
port 97 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 o_mem_write_M
port 98 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 o_pc_IF[0]
port 99 nsew signal output
rlabel metal3 s 79242 5448 80042 5568 6 o_pc_IF[10]
port 100 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 o_pc_IF[11]
port 101 nsew signal output
rlabel metal2 s 23846 78618 23902 79418 6 o_pc_IF[12]
port 102 nsew signal output
rlabel metal3 s 79242 40128 80042 40248 6 o_pc_IF[13]
port 103 nsew signal output
rlabel metal2 s 65706 78618 65762 79418 6 o_pc_IF[14]
port 104 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 o_pc_IF[15]
port 105 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 o_pc_IF[16]
port 106 nsew signal output
rlabel metal3 s 79242 42168 80042 42288 6 o_pc_IF[17]
port 107 nsew signal output
rlabel metal2 s 33506 78618 33562 79418 6 o_pc_IF[18]
port 108 nsew signal output
rlabel metal3 s 79242 27888 80042 28008 6 o_pc_IF[19]
port 109 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 o_pc_IF[1]
port 110 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 o_pc_IF[20]
port 111 nsew signal output
rlabel metal3 s 79242 53728 80042 53848 6 o_pc_IF[21]
port 112 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 o_pc_IF[22]
port 113 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 o_pc_IF[23]
port 114 nsew signal output
rlabel metal3 s 79242 19728 80042 19848 6 o_pc_IF[24]
port 115 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 o_pc_IF[25]
port 116 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 o_pc_IF[26]
port 117 nsew signal output
rlabel metal2 s 18050 78618 18106 79418 6 o_pc_IF[27]
port 118 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 o_pc_IF[28]
port 119 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 o_pc_IF[29]
port 120 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 o_pc_IF[2]
port 121 nsew signal output
rlabel metal3 s 79242 11568 80042 11688 6 o_pc_IF[30]
port 122 nsew signal output
rlabel metal3 s 79242 65968 80042 66088 6 o_pc_IF[31]
port 123 nsew signal output
rlabel metal3 s 79242 46248 80042 46368 6 o_pc_IF[3]
port 124 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 o_pc_IF[4]
port 125 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 o_pc_IF[5]
port 126 nsew signal output
rlabel metal3 s 79242 23808 80042 23928 6 o_pc_IF[6]
port 127 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 o_pc_IF[7]
port 128 nsew signal output
rlabel metal3 s 79242 49648 80042 49768 6 o_pc_IF[8]
port 129 nsew signal output
rlabel metal3 s 79242 74128 80042 74248 6 o_pc_IF[9]
port 130 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 o_write_data_M[0]
port 131 nsew signal output
rlabel metal3 s 79242 78208 80042 78328 6 o_write_data_M[10]
port 132 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 o_write_data_M[11]
port 133 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 o_write_data_M[12]
port 134 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 o_write_data_M[13]
port 135 nsew signal output
rlabel metal2 s 18 0 74 800 6 o_write_data_M[14]
port 136 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 o_write_data_M[15]
port 137 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 o_write_data_M[16]
port 138 nsew signal output
rlabel metal2 s 16118 78618 16174 79418 6 o_write_data_M[17]
port 139 nsew signal output
rlabel metal2 s 43166 78618 43222 79418 6 o_write_data_M[18]
port 140 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 o_write_data_M[19]
port 141 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 o_write_data_M[1]
port 142 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 o_write_data_M[20]
port 143 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 o_write_data_M[21]
port 144 nsew signal output
rlabel metal2 s 41234 78618 41290 79418 6 o_write_data_M[22]
port 145 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 o_write_data_M[23]
port 146 nsew signal output
rlabel metal2 s 67638 78618 67694 79418 6 o_write_data_M[24]
port 147 nsew signal output
rlabel metal3 s 79242 13608 80042 13728 6 o_write_data_M[25]
port 148 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 o_write_data_M[26]
port 149 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 o_write_data_M[27]
port 150 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 o_write_data_M[28]
port 151 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 o_write_data_M[29]
port 152 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 o_write_data_M[2]
port 153 nsew signal output
rlabel metal3 s 79242 51688 80042 51808 6 o_write_data_M[30]
port 154 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 o_write_data_M[31]
port 155 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 o_write_data_M[3]
port 156 nsew signal output
rlabel metal2 s 57978 78618 58034 79418 6 o_write_data_M[4]
port 157 nsew signal output
rlabel metal2 s 662 78618 718 79418 6 o_write_data_M[5]
port 158 nsew signal output
rlabel metal2 s 14186 78618 14242 79418 6 o_write_data_M[6]
port 159 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 o_write_data_M[7]
port 160 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 o_write_data_M[8]
port 161 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 o_write_data_M[9]
port 162 nsew signal output
rlabel metal3 s 79242 38088 80042 38208 6 rst
port 163 nsew signal input
rlabel metal4 s 5864 2672 6184 76752 6 vccd1
port 164 nsew power bidirectional
rlabel metal4 s 36584 2672 36904 76752 6 vccd1
port 164 nsew power bidirectional
rlabel metal4 s 67304 2672 67624 76752 6 vccd1
port 164 nsew power bidirectional
rlabel metal4 s 6524 2672 6844 76752 6 vssd1
port 165 nsew ground bidirectional
rlabel metal4 s 37244 2672 37564 76752 6 vssd1
port 165 nsew ground bidirectional
rlabel metal4 s 67964 2672 68284 76752 6 vssd1
port 165 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 80042 79418
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 23034502
string GDS_FILE /home/roliveira/Desktop/osiris_i/openlane/core/runs/metal/results/signoff/core.magic.gds
string GDS_START 923568
<< end >>

