// This is the unpowered netlist.
module uart_wbs_bridge (clk,
    i_start_rx,
    i_uart_rx,
    o_uart_tx,
    rst,
    wb_ack_i,
    wb_cyc_o,
    wb_stb_o,
    wb_we_o,
    wb_adr_o,
    wb_dat_i,
    wb_dat_o);
 input clk;
 input i_start_rx;
 input i_uart_rx;
 output o_uart_tx;
 input rst;
 input wb_ack_i;
 output wb_cyc_o;
 output wb_stb_o;
 output wb_we_o;
 output [31:0] wb_adr_o;
 input [31:0] wb_dat_i;
 output [31:0] wb_dat_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire \addr_reg[0] ;
 wire \addr_reg[10] ;
 wire \addr_reg[11] ;
 wire \addr_reg[12] ;
 wire \addr_reg[13] ;
 wire \addr_reg[14] ;
 wire \addr_reg[15] ;
 wire \addr_reg[16] ;
 wire \addr_reg[17] ;
 wire \addr_reg[18] ;
 wire \addr_reg[19] ;
 wire \addr_reg[1] ;
 wire \addr_reg[20] ;
 wire \addr_reg[21] ;
 wire \addr_reg[22] ;
 wire \addr_reg[23] ;
 wire \addr_reg[24] ;
 wire \addr_reg[25] ;
 wire \addr_reg[26] ;
 wire \addr_reg[27] ;
 wire \addr_reg[28] ;
 wire \addr_reg[29] ;
 wire \addr_reg[2] ;
 wire \addr_reg[30] ;
 wire \addr_reg[31] ;
 wire \addr_reg[3] ;
 wire \addr_reg[4] ;
 wire \addr_reg[5] ;
 wire \addr_reg[6] ;
 wire \addr_reg[7] ;
 wire \addr_reg[8] ;
 wire \addr_reg[9] ;
 wire \byte_count[0] ;
 wire \byte_count[1] ;
 wire \byte_count[2] ;
 wire \byte_count[3] ;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \cmd_reg[0] ;
 wire \cmd_reg[1] ;
 wire \cmd_reg[2] ;
 wire \cmd_reg[3] ;
 wire \cmd_reg[4] ;
 wire \cmd_reg[5] ;
 wire \cmd_reg[6] ;
 wire \cmd_reg[7] ;
 wire \data_reg[0] ;
 wire \data_reg[10] ;
 wire \data_reg[11] ;
 wire \data_reg[12] ;
 wire \data_reg[13] ;
 wire \data_reg[14] ;
 wire \data_reg[15] ;
 wire \data_reg[16] ;
 wire \data_reg[17] ;
 wire \data_reg[18] ;
 wire \data_reg[19] ;
 wire \data_reg[1] ;
 wire \data_reg[20] ;
 wire \data_reg[21] ;
 wire \data_reg[22] ;
 wire \data_reg[23] ;
 wire \data_reg[2] ;
 wire \data_reg[3] ;
 wire \data_reg[4] ;
 wire \data_reg[5] ;
 wire \data_reg[6] ;
 wire \data_reg[7] ;
 wire \data_reg[8] ;
 wire \data_reg[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \uart_rx_inst.bit_index[0] ;
 wire \uart_rx_inst.bit_index[1] ;
 wire \uart_rx_inst.bit_index[2] ;
 wire \uart_rx_inst.bit_index[3] ;
 wire \uart_rx_inst.clock_count[0] ;
 wire \uart_rx_inst.clock_count[10] ;
 wire \uart_rx_inst.clock_count[11] ;
 wire \uart_rx_inst.clock_count[12] ;
 wire \uart_rx_inst.clock_count[13] ;
 wire \uart_rx_inst.clock_count[14] ;
 wire \uart_rx_inst.clock_count[15] ;
 wire \uart_rx_inst.clock_count[1] ;
 wire \uart_rx_inst.clock_count[2] ;
 wire \uart_rx_inst.clock_count[3] ;
 wire \uart_rx_inst.clock_count[4] ;
 wire \uart_rx_inst.clock_count[5] ;
 wire \uart_rx_inst.clock_count[6] ;
 wire \uart_rx_inst.clock_count[7] ;
 wire \uart_rx_inst.clock_count[8] ;
 wire \uart_rx_inst.clock_count[9] ;
 wire \uart_rx_inst.o_data[0] ;
 wire \uart_rx_inst.o_data[1] ;
 wire \uart_rx_inst.o_data[2] ;
 wire \uart_rx_inst.o_data[3] ;
 wire \uart_rx_inst.o_data[4] ;
 wire \uart_rx_inst.o_data[5] ;
 wire \uart_rx_inst.o_data[6] ;
 wire \uart_rx_inst.o_data[7] ;
 wire \uart_rx_inst.o_data_valid ;
 wire \uart_rx_inst.receiving ;
 wire \uart_rx_inst.rx_sync_1 ;
 wire \uart_rx_inst.rx_sync_2 ;
 wire \uart_rx_inst.shift_reg[0] ;
 wire \uart_rx_inst.shift_reg[1] ;
 wire \uart_rx_inst.shift_reg[2] ;
 wire \uart_rx_inst.shift_reg[3] ;
 wire \uart_rx_inst.shift_reg[4] ;
 wire \uart_rx_inst.shift_reg[5] ;
 wire \uart_rx_inst.shift_reg[6] ;
 wire \uart_rx_inst.shift_reg[7] ;
 wire \uart_tx_inst.bit_index[0] ;
 wire \uart_tx_inst.bit_index[1] ;
 wire \uart_tx_inst.bit_index[2] ;
 wire \uart_tx_inst.bit_index[3] ;
 wire \uart_tx_inst.clock_count[0] ;
 wire \uart_tx_inst.clock_count[10] ;
 wire \uart_tx_inst.clock_count[11] ;
 wire \uart_tx_inst.clock_count[12] ;
 wire \uart_tx_inst.clock_count[13] ;
 wire \uart_tx_inst.clock_count[14] ;
 wire \uart_tx_inst.clock_count[15] ;
 wire \uart_tx_inst.clock_count[1] ;
 wire \uart_tx_inst.clock_count[2] ;
 wire \uart_tx_inst.clock_count[3] ;
 wire \uart_tx_inst.clock_count[4] ;
 wire \uart_tx_inst.clock_count[5] ;
 wire \uart_tx_inst.clock_count[6] ;
 wire \uart_tx_inst.clock_count[7] ;
 wire \uart_tx_inst.clock_count[8] ;
 wire \uart_tx_inst.clock_count[9] ;
 wire \uart_tx_inst.i_data[0] ;
 wire \uart_tx_inst.i_data[1] ;
 wire \uart_tx_inst.i_data[2] ;
 wire \uart_tx_inst.i_data[3] ;
 wire \uart_tx_inst.i_data[4] ;
 wire \uart_tx_inst.i_data[5] ;
 wire \uart_tx_inst.i_data[6] ;
 wire \uart_tx_inst.i_data[7] ;
 wire \uart_tx_inst.i_data_valid ;
 wire \uart_tx_inst.o_ready ;
 wire \uart_tx_inst.shift_reg[1] ;
 wire \uart_tx_inst.shift_reg[2] ;
 wire \uart_tx_inst.shift_reg[3] ;
 wire \uart_tx_inst.shift_reg[4] ;
 wire \uart_tx_inst.shift_reg[5] ;
 wire \uart_tx_inst.shift_reg[6] ;
 wire \uart_tx_inst.shift_reg[7] ;
 wire \uart_tx_inst.shift_reg[8] ;
 wire \uart_tx_inst.shift_reg[9] ;
 wire \uart_tx_inst.transmitting ;

 sky130_fd_sc_hd__diode_2 ANTENNA__0871__A0 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__A0 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__0948__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0948__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0949__C (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0955__A_N (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0956__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0957__A_N (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0957__C (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0957__D (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0962__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0962__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0964__A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0965__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__A0 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0969__C (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0971__C (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0972__A2_N (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0973__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0973__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0973__C_N (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__0974__A1_N (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0974__A2_N (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0974__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__C_N (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__0976__A1_N (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0976__A2_N (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0976__B2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0977__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0977__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__A1_N (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__B2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__C_N (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__A1_N (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__B2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__A1_N (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0983__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0983__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0983__C_N (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__A1_N (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__A1_N (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0989__A_N (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0989__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__A_N (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__C (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__0993__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__C (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__0997__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__A_N (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__A_N (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__C (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__1002__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__1003__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__1005__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__1006__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1006__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1006__B2 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1007__A_N (.DIODE(\byte_count[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1007__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__1007__C (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__A_N (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__1011__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1013__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1014__B1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__A (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__B1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__B2 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1017__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__1017__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1018__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1018__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1019__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1020__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1020__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1024__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1024__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1024__B2 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1025__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1026__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1026__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1027__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1028__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1028__B2 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__C (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__C (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__B2 (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__B2 (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1034__B2 (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__B2 (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1036__B2 (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__B2 (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__B2 (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__B2 (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1040__A2_N (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1041__A1_N (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1041__A2_N (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1041__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1042__A1_N (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1042__A2_N (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1042__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1043__A2_N (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1043__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1044__A2_N (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1044__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__A2_N (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1046__A2_N (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1046__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__A2_N (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1048__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1048__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1050__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1050__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1051__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1051__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1052__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1052__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1053__B1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1053__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1054__A1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__1054__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1054__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1055__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1055__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1056__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1056__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1057__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1057__B1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1057__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1058__B2 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1059__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1059__B2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__1060__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1060__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1061__B1 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1061__B2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__1062__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1063__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1063__B1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1063__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1064__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1065__A0 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__1065__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1066__A0 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__1066__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1067__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1068__A0 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__1069__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1070__A0 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__1070__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1071__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1075__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__1076__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1076__S0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__1076__S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1079__A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__1079__S0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__1079__S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__S0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1085__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1085__S0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__1085__S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__S0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__S0 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__S0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__S0 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__S1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1100__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__1100__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1100__C (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__1103__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1104__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__A0 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1106__A0 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__1106__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1107__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__A0 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1109__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__A0 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1111__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1112__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1115__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1116__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1118__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1120__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1121__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1122__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1124__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1125__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1126__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1127__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1128__S (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1129__S (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1130__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1131__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1132__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1133__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1134__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1135__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1142__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1143__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1145__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1146__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1156__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1158__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1160__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1161__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1164__A0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__1164__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1166__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1168__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__S (.DIODE(_0468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1170__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__S (.DIODE(_0468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1172__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__B1_N (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1178__A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__B1_N (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__1193__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__1194__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__1194__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__1340__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1416__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(_0468_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold115_A (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold165_A (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold173_A (.DIODE(\byte_count[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold204_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_95 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__inv_2 _0709_ (.A(net477),
    .Y(_0488_));
 sky130_fd_sc_hd__inv_2 _0710_ (.A(net278),
    .Y(_0489_));
 sky130_fd_sc_hd__inv_2 _0711_ (.A(net189),
    .Y(_0490_));
 sky130_fd_sc_hd__inv_2 _0712_ (.A(net325),
    .Y(_0491_));
 sky130_fd_sc_hd__inv_2 _0713_ (.A(net429),
    .Y(_0492_));
 sky130_fd_sc_hd__inv_2 _0714_ (.A(net433),
    .Y(_0493_));
 sky130_fd_sc_hd__inv_2 _0715_ (.A(net469),
    .Y(_0494_));
 sky130_fd_sc_hd__inv_2 _0716_ (.A(net482),
    .Y(_0495_));
 sky130_fd_sc_hd__inv_2 _0717_ (.A(net442),
    .Y(_0496_));
 sky130_fd_sc_hd__inv_2 _0718_ (.A(net494),
    .Y(_0497_));
 sky130_fd_sc_hd__inv_2 _0719_ (.A(net312),
    .Y(_0498_));
 sky130_fd_sc_hd__inv_2 _0720_ (.A(net4),
    .Y(_0499_));
 sky130_fd_sc_hd__inv_2 _0721_ (.A(net396),
    .Y(_0500_));
 sky130_fd_sc_hd__inv_2 _0722_ (.A(net121),
    .Y(_0003_));
 sky130_fd_sc_hd__nor2_1 _0723_ (.A(net325),
    .B(net429),
    .Y(_0501_));
 sky130_fd_sc_hd__or2_2 _0724_ (.A(net325),
    .B(net429),
    .X(_0502_));
 sky130_fd_sc_hd__or2_1 _0725_ (.A(net332),
    .B(net189),
    .X(_0503_));
 sky130_fd_sc_hd__nor2_1 _0726_ (.A(_0502_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__o21a_1 _0727_ (.A1(net189),
    .A2(_0502_),
    .B1(net332),
    .X(_0505_));
 sky130_fd_sc_hd__inv_2 _0728_ (.A(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__or4b_1 _0729_ (.A(net382),
    .B(net380),
    .C(net469),
    .D_N(net436),
    .X(_0507_));
 sky130_fd_sc_hd__or4bb_1 _0730_ (.A(net433),
    .B(\uart_rx_inst.clock_count[14] ),
    .C_N(\uart_rx_inst.clock_count[2] ),
    .D_N(\uart_rx_inst.clock_count[0] ),
    .X(_0508_));
 sky130_fd_sc_hd__or4_1 _0731_ (.A(net402),
    .B(\uart_rx_inst.clock_count[4] ),
    .C(net483),
    .D(\uart_rx_inst.clock_count[1] ),
    .X(_0509_));
 sky130_fd_sc_hd__or4b_1 _0732_ (.A(net424),
    .B(net416),
    .C(net479),
    .D_N(\uart_rx_inst.clock_count[6] ),
    .X(_0510_));
 sky130_fd_sc_hd__or4_1 _0733_ (.A(_0507_),
    .B(net434),
    .C(net484),
    .D(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__or2_2 _0734_ (.A(_0500_),
    .B(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__nor2_1 _0735_ (.A(_0505_),
    .B(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__or4_4 _0736_ (.A(_0500_),
    .B(_0504_),
    .C(_0505_),
    .D(net435),
    .X(_0514_));
 sky130_fd_sc_hd__or4_1 _0737_ (.A(net424),
    .B(net416),
    .C(net402),
    .D(net496),
    .X(_0515_));
 sky130_fd_sc_hd__or4bb_1 _0738_ (.A(net442),
    .B(net463),
    .C_N(\uart_rx_inst.clock_count[0] ),
    .D_N(net438),
    .X(_0516_));
 sky130_fd_sc_hd__or4b_1 _0739_ (.A(net433),
    .B(net450),
    .C(net479),
    .D_N(net458),
    .X(_0517_));
 sky130_fd_sc_hd__or4_1 _0740_ (.A(_0507_),
    .B(_0515_),
    .C(_0516_),
    .D(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__or4_1 _0741_ (.A(_0500_),
    .B(_0504_),
    .C(_0505_),
    .D(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__o31a_1 _0742_ (.A1(net189),
    .A2(_0502_),
    .A3(_0514_),
    .B1(net274),
    .X(_0520_));
 sky130_fd_sc_hd__xnor2_1 _0743_ (.A(net189),
    .B(net325),
    .Y(_0521_));
 sky130_fd_sc_hd__o21a_1 _0744_ (.A1(_0502_),
    .A2(_0503_),
    .B1(net165),
    .X(_0522_));
 sky130_fd_sc_hd__and2b_1 _0745_ (.A_N(_0519_),
    .B(_0521_),
    .X(_0523_));
 sky130_fd_sc_hd__a31o_1 _0746_ (.A1(net165),
    .A2(_0501_),
    .A3(_0523_),
    .B1(_0520_),
    .X(_0433_));
 sky130_fd_sc_hd__nand2_1 _0747_ (.A(net325),
    .B(net429),
    .Y(_0524_));
 sky130_fd_sc_hd__or2_1 _0748_ (.A(_0490_),
    .B(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__nor2_1 _0749_ (.A(_0514_),
    .B(net190),
    .Y(_0526_));
 sky130_fd_sc_hd__mux2_1 _0750_ (.A0(net139),
    .A1(net165),
    .S(net191),
    .X(_0432_));
 sky130_fd_sc_hd__and4bb_1 _0751_ (.A_N(\uart_rx_inst.bit_index[0] ),
    .B_N(_0514_),
    .C(\uart_rx_inst.bit_index[2] ),
    .D(\uart_rx_inst.bit_index[1] ),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _0752_ (.A0(net137),
    .A1(net165),
    .S(_0527_),
    .X(_0431_));
 sky130_fd_sc_hd__or4_1 _0753_ (.A(_0490_),
    .B(\uart_rx_inst.bit_index[1] ),
    .C(_0492_),
    .D(_0514_),
    .X(_0528_));
 sky130_fd_sc_hd__and4_1 _0754_ (.A(_0491_),
    .B(\uart_rx_inst.bit_index[0] ),
    .C(\uart_rx_inst.rx_sync_2 ),
    .D(_0503_),
    .X(_0529_));
 sky130_fd_sc_hd__and2b_1 _0755_ (.A_N(_0514_),
    .B(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__a21o_1 _0756_ (.A1(net159),
    .A2(_0528_),
    .B1(_0530_),
    .X(_0430_));
 sky130_fd_sc_hd__o31a_1 _0757_ (.A1(_0490_),
    .A2(_0502_),
    .A3(_0514_),
    .B1(net343),
    .X(_0531_));
 sky130_fd_sc_hd__nor2_1 _0758_ (.A(_0519_),
    .B(_0521_),
    .Y(_0532_));
 sky130_fd_sc_hd__a31o_1 _0759_ (.A1(_0501_),
    .A2(_0522_),
    .A3(_0532_),
    .B1(_0531_),
    .X(_0429_));
 sky130_fd_sc_hd__o31a_1 _0760_ (.A1(_0503_),
    .A2(_0514_),
    .A3(_0524_),
    .B1(net151),
    .X(_0533_));
 sky130_fd_sc_hd__a41o_1 _0761_ (.A1(net325),
    .A2(net429),
    .A3(net165),
    .A4(_0532_),
    .B1(_0533_),
    .X(_0428_));
 sky130_fd_sc_hd__o41a_1 _0762_ (.A1(_0491_),
    .A2(net429),
    .A3(_0514_),
    .A4(_0521_),
    .B1(net345),
    .X(_0534_));
 sky130_fd_sc_hd__a41o_1 _0763_ (.A1(net325),
    .A2(_0492_),
    .A3(net165),
    .A4(_0532_),
    .B1(_0534_),
    .X(_0427_));
 sky130_fd_sc_hd__or4_1 _0764_ (.A(net325),
    .B(_0492_),
    .C(_0503_),
    .D(_0519_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _0765_ (.A0(_0522_),
    .A1(net175),
    .S(net326),
    .X(_0426_));
 sky130_fd_sc_hd__and2_1 _0766_ (.A(net426),
    .B(\uart_tx_inst.bit_index[0] ),
    .X(_0536_));
 sky130_fd_sc_hd__nand2_1 _0767_ (.A(net426),
    .B(net452),
    .Y(_0537_));
 sky130_fd_sc_hd__nand2_1 _0768_ (.A(net413),
    .B(net427),
    .Y(_0538_));
 sky130_fd_sc_hd__or4b_1 _0769_ (.A(net446),
    .B(net362),
    .C(net409),
    .D_N(net431),
    .X(_0539_));
 sky130_fd_sc_hd__or4bb_1 _0770_ (.A(\uart_tx_inst.clock_count[15] ),
    .B(\uart_tx_inst.clock_count[14] ),
    .C_N(net419),
    .D_N(\uart_tx_inst.clock_count[0] ),
    .X(_0540_));
 sky130_fd_sc_hd__or4_1 _0771_ (.A(\uart_tx_inst.clock_count[5] ),
    .B(\uart_tx_inst.clock_count[4] ),
    .C(net405),
    .D(\uart_tx_inst.clock_count[1] ),
    .X(_0541_));
 sky130_fd_sc_hd__or4b_1 _0772_ (.A(\uart_tx_inst.clock_count[9] ),
    .B(\uart_tx_inst.clock_count[8] ),
    .C(\uart_tx_inst.clock_count[7] ),
    .D_N(net444),
    .X(_0542_));
 sky130_fd_sc_hd__or4_1 _0773_ (.A(_0539_),
    .B(_0540_),
    .C(_0541_),
    .D(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__nor2_2 _0774_ (.A(_0497_),
    .B(net447),
    .Y(_0544_));
 sky130_fd_sc_hd__nand2_1 _0775_ (.A(net391),
    .B(net241),
    .Y(_0545_));
 sky130_fd_sc_hd__and2_2 _0776_ (.A(_0497_),
    .B(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__or4b_1 _0777_ (.A(net475),
    .B(net495),
    .C(net454),
    .D_N(net444),
    .X(_0547_));
 sky130_fd_sc_hd__or4bb_1 _0778_ (.A(net405),
    .B(net456),
    .C_N(\uart_tx_inst.clock_count[0] ),
    .D_N(net419),
    .X(_0548_));
 sky130_fd_sc_hd__or4_1 _0779_ (.A(net362),
    .B(net409),
    .C(net472),
    .D(net491),
    .X(_0549_));
 sky130_fd_sc_hd__or4b_1 _0780_ (.A(net477),
    .B(net487),
    .C(net446),
    .D_N(net431),
    .X(_0550_));
 sky130_fd_sc_hd__or4_1 _0781_ (.A(_0547_),
    .B(_0548_),
    .C(_0549_),
    .D(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__and2_1 _0782_ (.A(\uart_tx_inst.transmitting ),
    .B(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__a21o_1 _0783_ (.A1(net494),
    .A2(_0551_),
    .B1(_0546_),
    .X(_0553_));
 sky130_fd_sc_hd__and2_1 _0784_ (.A(_0538_),
    .B(_0544_),
    .X(_0554_));
 sky130_fd_sc_hd__a21o_1 _0785_ (.A1(_0538_),
    .A2(_0544_),
    .B1(_0553_),
    .X(_0555_));
 sky130_fd_sc_hd__nor2_1 _0786_ (.A(net356),
    .B(_0538_),
    .Y(_0556_));
 sky130_fd_sc_hd__a22o_1 _0787_ (.A1(net356),
    .A2(_0555_),
    .B1(_0556_),
    .B2(net448),
    .X(_0425_));
 sky130_fd_sc_hd__a22o_1 _0788_ (.A1(net427),
    .A2(_0554_),
    .B1(_0555_),
    .B2(net413),
    .X(_0424_));
 sky130_fd_sc_hd__or2_1 _0789_ (.A(net426),
    .B(net452),
    .X(_0557_));
 sky130_fd_sc_hd__a32o_1 _0790_ (.A1(_0537_),
    .A2(net448),
    .A3(_0557_),
    .B1(_0553_),
    .B2(net426),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _0791_ (.A0(_0553_),
    .A1(net448),
    .S(net452),
    .X(_0558_));
 sky130_fd_sc_hd__inv_2 _0792_ (.A(_0558_),
    .Y(_0422_));
 sky130_fd_sc_hd__nand2_1 _0793_ (.A(net456),
    .B(\uart_tx_inst.clock_count[0] ),
    .Y(_0559_));
 sky130_fd_sc_hd__nand3_1 _0794_ (.A(net419),
    .B(\uart_tx_inst.clock_count[1] ),
    .C(\uart_tx_inst.clock_count[0] ),
    .Y(_0560_));
 sky130_fd_sc_hd__and4_2 _0795_ (.A(net405),
    .B(net419),
    .C(net456),
    .D(net485),
    .X(_0561_));
 sky130_fd_sc_hd__inv_2 _0796_ (.A(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__nand2_1 _0797_ (.A(net454),
    .B(_0561_),
    .Y(_0563_));
 sky130_fd_sc_hd__and3_1 _0798_ (.A(net475),
    .B(net444),
    .C(net497),
    .X(_0564_));
 sky130_fd_sc_hd__and4_1 _0799_ (.A(net491),
    .B(net454),
    .C(_0561_),
    .D(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__nor2_4 _0800_ (.A(\uart_tx_inst.transmitting ),
    .B(_0545_),
    .Y(_0566_));
 sky130_fd_sc_hd__or2_2 _0801_ (.A(net494),
    .B(_0545_),
    .X(_0567_));
 sky130_fd_sc_hd__nor2_1 _0802_ (.A(_0488_),
    .B(_0566_),
    .Y(_0568_));
 sky130_fd_sc_hd__and4_1 _0803_ (.A(net362),
    .B(net409),
    .C(net472),
    .D(net491),
    .X(_0569_));
 sky130_fd_sc_hd__and4_1 _0804_ (.A(net454),
    .B(_0561_),
    .C(_0564_),
    .D(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__nand2_1 _0805_ (.A(net431),
    .B(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__and4_1 _0806_ (.A(net446),
    .B(net431),
    .C(net494),
    .D(_0570_),
    .X(_0572_));
 sky130_fd_sc_hd__nand2_1 _0807_ (.A(net487),
    .B(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__mux2_1 _0808_ (.A0(_0488_),
    .A1(_0568_),
    .S(_0573_),
    .X(_0421_));
 sky130_fd_sc_hd__o21a_1 _0809_ (.A1(net487),
    .A2(_0572_),
    .B1(_0567_),
    .X(_0574_));
 sky130_fd_sc_hd__and2_1 _0810_ (.A(net488),
    .B(_0574_),
    .X(_0420_));
 sky130_fd_sc_hd__o2bb2a_1 _0811_ (.A1_N(net446),
    .A2_N(_0567_),
    .B1(_0571_),
    .B2(_0497_),
    .X(_0575_));
 sky130_fd_sc_hd__nor2_1 _0812_ (.A(_0572_),
    .B(_0575_),
    .Y(_0419_));
 sky130_fd_sc_hd__or2_1 _0813_ (.A(net431),
    .B(_0570_),
    .X(_0576_));
 sky130_fd_sc_hd__a32o_1 _0814_ (.A1(_0552_),
    .A2(_0571_),
    .A3(_0576_),
    .B1(_0546_),
    .B2(net431),
    .X(_0418_));
 sky130_fd_sc_hd__nand2_1 _0815_ (.A(\uart_tx_inst.transmitting ),
    .B(_0565_),
    .Y(_0577_));
 sky130_fd_sc_hd__and3_1 _0816_ (.A(net472),
    .B(\uart_tx_inst.transmitting ),
    .C(_0565_),
    .X(_0578_));
 sky130_fd_sc_hd__and4_1 _0817_ (.A(net409),
    .B(\uart_tx_inst.clock_count[9] ),
    .C(\uart_tx_inst.transmitting ),
    .D(_0565_),
    .X(_0579_));
 sky130_fd_sc_hd__o21ai_1 _0818_ (.A1(net362),
    .A2(_0579_),
    .B1(_0567_),
    .Y(_0580_));
 sky130_fd_sc_hd__a21oi_1 _0819_ (.A1(net362),
    .A2(_0579_),
    .B1(_0580_),
    .Y(_0417_));
 sky130_fd_sc_hd__nor2_1 _0820_ (.A(_0566_),
    .B(_0579_),
    .Y(_0581_));
 sky130_fd_sc_hd__o21a_1 _0821_ (.A1(net409),
    .A2(_0578_),
    .B1(_0581_),
    .X(_0416_));
 sky130_fd_sc_hd__nand2_1 _0822_ (.A(net472),
    .B(_0567_),
    .Y(_0582_));
 sky130_fd_sc_hd__a21oi_1 _0823_ (.A1(_0577_),
    .A2(net473),
    .B1(_0578_),
    .Y(_0415_));
 sky130_fd_sc_hd__a41o_1 _0824_ (.A1(net454),
    .A2(\uart_tx_inst.transmitting ),
    .A3(_0561_),
    .A4(_0564_),
    .B1(net491),
    .X(_0583_));
 sky130_fd_sc_hd__and3_1 _0825_ (.A(_0567_),
    .B(_0577_),
    .C(net492),
    .X(_0414_));
 sky130_fd_sc_hd__and3_1 _0826_ (.A(net454),
    .B(net494),
    .C(_0561_),
    .X(_0584_));
 sky130_fd_sc_hd__and3_1 _0827_ (.A(net444),
    .B(\uart_tx_inst.clock_count[5] ),
    .C(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__nand2_1 _0828_ (.A(net475),
    .B(_0567_),
    .Y(_0586_));
 sky130_fd_sc_hd__mux2_1 _0829_ (.A0(_0586_),
    .A1(net475),
    .S(_0585_),
    .X(_0587_));
 sky130_fd_sc_hd__inv_2 _0830_ (.A(net476),
    .Y(_0413_));
 sky130_fd_sc_hd__or3b_1 _0831_ (.A(_0546_),
    .B(_0563_),
    .C_N(\uart_tx_inst.clock_count[5] ),
    .X(_0588_));
 sky130_fd_sc_hd__nand2_1 _0832_ (.A(net495),
    .B(_0584_),
    .Y(_0589_));
 sky130_fd_sc_hd__nor2_1 _0833_ (.A(net444),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__a31o_1 _0834_ (.A1(net444),
    .A2(_0553_),
    .A3(_0588_),
    .B1(_0590_),
    .X(_0412_));
 sky130_fd_sc_hd__or2_1 _0835_ (.A(net495),
    .B(_0584_),
    .X(_0591_));
 sky130_fd_sc_hd__and3_1 _0836_ (.A(_0567_),
    .B(_0589_),
    .C(_0591_),
    .X(_0411_));
 sky130_fd_sc_hd__or2_1 _0837_ (.A(net454),
    .B(_0561_),
    .X(_0592_));
 sky130_fd_sc_hd__a32o_1 _0838_ (.A1(\uart_tx_inst.transmitting ),
    .A2(_0563_),
    .A3(_0592_),
    .B1(_0546_),
    .B2(net454),
    .X(_0410_));
 sky130_fd_sc_hd__a31o_1 _0839_ (.A1(\uart_tx_inst.clock_count[2] ),
    .A2(\uart_tx_inst.clock_count[1] ),
    .A3(\uart_tx_inst.clock_count[0] ),
    .B1(net405),
    .X(_0593_));
 sky130_fd_sc_hd__a32o_1 _0840_ (.A1(\uart_tx_inst.transmitting ),
    .A2(_0562_),
    .A3(_0593_),
    .B1(_0546_),
    .B2(net405),
    .X(_0409_));
 sky130_fd_sc_hd__a21o_1 _0841_ (.A1(\uart_tx_inst.clock_count[1] ),
    .A2(\uart_tx_inst.clock_count[0] ),
    .B1(net419),
    .X(_0594_));
 sky130_fd_sc_hd__a32o_1 _0842_ (.A1(_0552_),
    .A2(_0560_),
    .A3(_0594_),
    .B1(_0546_),
    .B2(net419),
    .X(_0408_));
 sky130_fd_sc_hd__or2_1 _0843_ (.A(net456),
    .B(\uart_tx_inst.clock_count[0] ),
    .X(_0595_));
 sky130_fd_sc_hd__a32o_1 _0844_ (.A1(_0552_),
    .A2(_0559_),
    .A3(_0595_),
    .B1(_0546_),
    .B2(net456),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _0845_ (.A0(\uart_tx_inst.transmitting ),
    .A1(_0546_),
    .S(net485),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _0846_ (.A0(net167),
    .A1(net259),
    .S(net452),
    .X(_0596_));
 sky130_fd_sc_hd__nor2_1 _0847_ (.A(net356),
    .B(net413),
    .Y(_0597_));
 sky130_fd_sc_hd__a32o_1 _0848_ (.A1(net452),
    .A2(\uart_tx_inst.shift_reg[1] ),
    .A3(_0597_),
    .B1(_0596_),
    .B2(net413),
    .X(_0598_));
 sky130_fd_sc_hd__and2b_1 _0849_ (.A_N(net426),
    .B(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__or2_1 _0850_ (.A(net413),
    .B(\uart_tx_inst.bit_index[1] ),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _0851_ (.A0(\uart_tx_inst.shift_reg[8] ),
    .A1(net147),
    .S(net452),
    .X(_0601_));
 sky130_fd_sc_hd__or2_1 _0852_ (.A(net414),
    .B(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__mux4_1 _0853_ (.A0(net183),
    .A1(\uart_tx_inst.shift_reg[3] ),
    .A2(net197),
    .A3(\uart_tx_inst.shift_reg[7] ),
    .S0(net452),
    .S1(net413),
    .X(_0603_));
 sky130_fd_sc_hd__a22o_1 _0854_ (.A1(net356),
    .A2(_0602_),
    .B1(_0603_),
    .B2(net426),
    .X(_0604_));
 sky130_fd_sc_hd__or2_1 _0855_ (.A(_0599_),
    .B(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__a22o_1 _0856_ (.A1(net466),
    .A2(_0553_),
    .B1(_0605_),
    .B2(net448),
    .X(_0405_));
 sky130_fd_sc_hd__or2_1 _0857_ (.A(net147),
    .B(_0566_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _0858_ (.A0(net500),
    .A1(net149),
    .S(_0566_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _0859_ (.A0(net501),
    .A1(net155),
    .S(_0566_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _0860_ (.A0(net197),
    .A1(net239),
    .S(_0566_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _0861_ (.A0(net259),
    .A1(net276),
    .S(_0566_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _0862_ (.A0(net167),
    .A1(net349),
    .S(_0566_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _0863_ (.A0(net503),
    .A1(net270),
    .S(_0566_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _0864_ (.A0(net183),
    .A1(net195),
    .S(_0566_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _0865_ (.A0(net504),
    .A1(net143),
    .S(_0566_),
    .X(_0396_));
 sky130_fd_sc_hd__nor2_4 _0866_ (.A(_0506_),
    .B(_0512_),
    .Y(_0000_));
 sky130_fd_sc_hd__mux2_1 _0867_ (.A0(net502),
    .A1(net274),
    .S(_0000_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _0868_ (.A0(\uart_rx_inst.o_data[6] ),
    .A1(net139),
    .S(_0000_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _0869_ (.A0(\uart_rx_inst.o_data[5] ),
    .A1(net137),
    .S(_0000_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _0870_ (.A0(net263),
    .A1(net159),
    .S(_0000_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _0871_ (.A0(net219),
    .A1(net343),
    .S(_0000_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _0872_ (.A0(net507),
    .A1(net151),
    .S(_0000_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _0873_ (.A0(net256),
    .A1(net345),
    .S(_0000_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _0874_ (.A0(net505),
    .A1(net175),
    .S(_0000_),
    .X(_0388_));
 sky130_fd_sc_hd__nand2_1 _0875_ (.A(net1),
    .B(_0500_),
    .Y(_0606_));
 sky130_fd_sc_hd__inv_2 _0876_ (.A(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__o31a_1 _0877_ (.A1(_0500_),
    .A2(_0505_),
    .A3(net480),
    .B1(_0606_),
    .X(_0608_));
 sky130_fd_sc_hd__a21o_1 _0878_ (.A1(net396),
    .A2(net190),
    .B1(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__a21o_1 _0879_ (.A1(net332),
    .A2(net397),
    .B1(net191),
    .X(_0387_));
 sky130_fd_sc_hd__nor2_1 _0880_ (.A(_0524_),
    .B(_0608_),
    .Y(_0610_));
 sky130_fd_sc_hd__o21a_1 _0881_ (.A1(net189),
    .A2(_0610_),
    .B1(net397),
    .X(_0386_));
 sky130_fd_sc_hd__or4b_1 _0882_ (.A(net332),
    .B(_0501_),
    .C(_0512_),
    .D_N(_0524_),
    .X(_0611_));
 sky130_fd_sc_hd__a21bo_1 _0883_ (.A1(net325),
    .A2(_0608_),
    .B1_N(_0611_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _0884_ (.A0(_0513_),
    .A1(_0608_),
    .S(net429),
    .X(_0384_));
 sky130_fd_sc_hd__nand3_1 _0885_ (.A(net438),
    .B(\uart_rx_inst.clock_count[1] ),
    .C(\uart_rx_inst.clock_count[0] ),
    .Y(_0612_));
 sky130_fd_sc_hd__and4_2 _0886_ (.A(net442),
    .B(net438),
    .C(net463),
    .D(net490),
    .X(_0613_));
 sky130_fd_sc_hd__and3_1 _0887_ (.A(net402),
    .B(net482),
    .C(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__inv_2 _0888_ (.A(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__and4_1 _0889_ (.A(\uart_rx_inst.clock_count[7] ),
    .B(net458),
    .C(net402),
    .D(\uart_rx_inst.clock_count[4] ),
    .X(_0616_));
 sky130_fd_sc_hd__and4_1 _0890_ (.A(net424),
    .B(net416),
    .C(_0613_),
    .D(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__nand2_1 _0891_ (.A(net469),
    .B(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__and3_2 _0892_ (.A(net380),
    .B(net469),
    .C(_0617_),
    .X(_0619_));
 sky130_fd_sc_hd__and2_1 _0893_ (.A(net382),
    .B(net436),
    .X(_0620_));
 sky130_fd_sc_hd__nand2_1 _0894_ (.A(_0619_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__nand3_1 _0895_ (.A(net450),
    .B(_0619_),
    .C(_0620_),
    .Y(_0622_));
 sky130_fd_sc_hd__and4_1 _0896_ (.A(net450),
    .B(net396),
    .C(_0619_),
    .D(_0620_),
    .X(_0623_));
 sky130_fd_sc_hd__nor2_1 _0897_ (.A(_0493_),
    .B(_0607_),
    .Y(_0624_));
 sky130_fd_sc_hd__mux2_1 _0898_ (.A0(_0624_),
    .A1(_0493_),
    .S(_0623_),
    .X(_0383_));
 sky130_fd_sc_hd__nor2_2 _0899_ (.A(net1),
    .B(net396),
    .Y(_0625_));
 sky130_fd_sc_hd__a21o_1 _0900_ (.A1(_0619_),
    .A2(_0620_),
    .B1(net450),
    .X(_0626_));
 sky130_fd_sc_hd__a32o_1 _0901_ (.A1(net396),
    .A2(_0622_),
    .A3(_0626_),
    .B1(_0625_),
    .B2(net450),
    .X(_0382_));
 sky130_fd_sc_hd__nand2_1 _0902_ (.A(net436),
    .B(_0619_),
    .Y(_0627_));
 sky130_fd_sc_hd__a21o_1 _0903_ (.A1(\uart_rx_inst.clock_count[12] ),
    .A2(_0619_),
    .B1(net382),
    .X(_0628_));
 sky130_fd_sc_hd__a32o_1 _0904_ (.A1(\uart_rx_inst.receiving ),
    .A2(_0621_),
    .A3(_0628_),
    .B1(_0625_),
    .B2(net382),
    .X(_0381_));
 sky130_fd_sc_hd__or2_1 _0905_ (.A(net436),
    .B(_0619_),
    .X(_0629_));
 sky130_fd_sc_hd__and2_1 _0906_ (.A(net396),
    .B(_0518_),
    .X(_0630_));
 sky130_fd_sc_hd__a32o_1 _0907_ (.A1(_0627_),
    .A2(_0629_),
    .A3(_0630_),
    .B1(_0625_),
    .B2(net436),
    .X(_0380_));
 sky130_fd_sc_hd__a21oi_1 _0908_ (.A1(net396),
    .A2(_0618_),
    .B1(_0625_),
    .Y(_0631_));
 sky130_fd_sc_hd__o2bb2a_1 _0909_ (.A1_N(\uart_rx_inst.receiving ),
    .A2_N(_0619_),
    .B1(_0631_),
    .B2(net380),
    .X(_0379_));
 sky130_fd_sc_hd__and3_1 _0910_ (.A(_0494_),
    .B(net396),
    .C(_0617_),
    .X(_0632_));
 sky130_fd_sc_hd__o21bai_1 _0911_ (.A1(_0494_),
    .A2(_0631_),
    .B1_N(_0632_),
    .Y(_0378_));
 sky130_fd_sc_hd__and4_1 _0912_ (.A(net416),
    .B(net396),
    .C(_0613_),
    .D(_0616_),
    .X(_0633_));
 sky130_fd_sc_hd__nor2_1 _0913_ (.A(_0607_),
    .B(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__mux2_1 _0914_ (.A0(_0633_),
    .A1(_0634_),
    .S(net424),
    .X(_0377_));
 sky130_fd_sc_hd__and4b_1 _0915_ (.A_N(net416),
    .B(net396),
    .C(_0613_),
    .D(_0616_),
    .X(_0635_));
 sky130_fd_sc_hd__a21o_1 _0916_ (.A1(net416),
    .A2(_0634_),
    .B1(_0635_),
    .X(_0376_));
 sky130_fd_sc_hd__nor2_1 _0917_ (.A(_0500_),
    .B(_0615_),
    .Y(_0636_));
 sky130_fd_sc_hd__and3_1 _0918_ (.A(net458),
    .B(net396),
    .C(_0614_),
    .X(_0637_));
 sky130_fd_sc_hd__nand2_1 _0919_ (.A(net479),
    .B(_0606_),
    .Y(_0638_));
 sky130_fd_sc_hd__mux2_1 _0920_ (.A0(_0638_),
    .A1(net479),
    .S(_0637_),
    .X(_0639_));
 sky130_fd_sc_hd__inv_2 _0921_ (.A(_0639_),
    .Y(_0375_));
 sky130_fd_sc_hd__a21o_1 _0922_ (.A1(_0615_),
    .A2(_0630_),
    .B1(_0625_),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _0923_ (.A0(_0636_),
    .A1(_0640_),
    .S(net458),
    .X(_0374_));
 sky130_fd_sc_hd__a21oi_1 _0924_ (.A1(net482),
    .A2(_0613_),
    .B1(_0500_),
    .Y(_0641_));
 sky130_fd_sc_hd__nor2_1 _0925_ (.A(_0625_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__o22a_1 _0926_ (.A1(_0500_),
    .A2(_0615_),
    .B1(_0642_),
    .B2(net402),
    .X(_0373_));
 sky130_fd_sc_hd__a2bb2o_1 _0927_ (.A1_N(_0495_),
    .A2_N(_0642_),
    .B1(_0641_),
    .B2(_0613_),
    .X(_0372_));
 sky130_fd_sc_hd__o2bb2a_1 _0928_ (.A1_N(net442),
    .A2_N(_0625_),
    .B1(_0613_),
    .B2(_0500_),
    .X(_0643_));
 sky130_fd_sc_hd__a21oi_1 _0929_ (.A1(_0496_),
    .A2(_0612_),
    .B1(_0643_),
    .Y(_0371_));
 sky130_fd_sc_hd__a21o_1 _0930_ (.A1(\uart_rx_inst.clock_count[1] ),
    .A2(\uart_rx_inst.clock_count[0] ),
    .B1(net438),
    .X(_0644_));
 sky130_fd_sc_hd__a32o_1 _0931_ (.A1(_0612_),
    .A2(_0630_),
    .A3(_0644_),
    .B1(_0625_),
    .B2(net438),
    .X(_0370_));
 sky130_fd_sc_hd__a21boi_1 _0932_ (.A1(net463),
    .A2(\uart_rx_inst.clock_count[0] ),
    .B1_N(_0518_),
    .Y(_0645_));
 sky130_fd_sc_hd__and2_1 _0933_ (.A(\uart_rx_inst.clock_count[0] ),
    .B(net396),
    .X(_0646_));
 sky130_fd_sc_hd__o32a_1 _0934_ (.A1(net463),
    .A2(_0607_),
    .A3(_0646_),
    .B1(_0645_),
    .B2(_0500_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _0935_ (.A0(_0625_),
    .A1(net396),
    .S(net490),
    .X(_0647_));
 sky130_fd_sc_hd__inv_2 _0936_ (.A(_0647_),
    .Y(_0368_));
 sky130_fd_sc_hd__and3b_2 _0937_ (.A_N(net481),
    .B(net312),
    .C(net411),
    .X(_0648_));
 sky130_fd_sc_hd__nand2b_1 _0938_ (.A_N(\uart_tx_inst.i_data_valid ),
    .B(net241),
    .Y(_0649_));
 sky130_fd_sc_hd__nand2b_1 _0939_ (.A_N(net312),
    .B(net411),
    .Y(_0650_));
 sky130_fd_sc_hd__a2bb2o_1 _0940_ (.A1_N(net4),
    .A2_N(_0650_),
    .B1(net242),
    .B2(_0648_),
    .X(_0651_));
 sky130_fd_sc_hd__and2b_1 _0941_ (.A_N(net312),
    .B(net418),
    .X(_0652_));
 sky130_fd_sc_hd__and3b_1 _0942_ (.A_N(net312),
    .B(net418),
    .C(net411),
    .X(_0653_));
 sky130_fd_sc_hd__and3b_1 _0943_ (.A_N(net411),
    .B(net312),
    .C(net418),
    .X(_0654_));
 sky130_fd_sc_hd__nor2_1 _0944_ (.A(net411),
    .B(net418),
    .Y(_0655_));
 sky130_fd_sc_hd__or4_1 _0945_ (.A(_0648_),
    .B(_0653_),
    .C(_0654_),
    .D(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__or3_1 _0946_ (.A(net411),
    .B(net299),
    .C(_0652_),
    .X(_0657_));
 sky130_fd_sc_hd__and3b_2 _0947_ (.A_N(_0651_),
    .B(_0656_),
    .C(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__nand2_1 _0948_ (.A(net116),
    .B(net118),
    .Y(_0659_));
 sky130_fd_sc_hd__and3_1 _0949_ (.A(net221),
    .B(net215),
    .C(net117),
    .X(_0660_));
 sky130_fd_sc_hd__nor3b_1 _0950_ (.A(net411),
    .B(net465),
    .C_N(net312),
    .Y(_0661_));
 sky130_fd_sc_hd__or3b_1 _0951_ (.A(\state[2] ),
    .B(\state[0] ),
    .C_N(net498),
    .X(_0662_));
 sky130_fd_sc_hd__or3_2 _0952_ (.A(_0648_),
    .B(_0654_),
    .C(_0661_),
    .X(_0663_));
 sky130_fd_sc_hd__inv_2 _0953_ (.A(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__o21ai_1 _0954_ (.A1(_0660_),
    .A2(_0664_),
    .B1(_0658_),
    .Y(_0665_));
 sky130_fd_sc_hd__and4b_1 _0955_ (.A_N(net115),
    .B(_0658_),
    .C(_0660_),
    .D(_0663_),
    .X(_0666_));
 sky130_fd_sc_hd__a21o_1 _0956_ (.A1(net115),
    .A2(_0665_),
    .B1(_0666_),
    .X(_0367_));
 sky130_fd_sc_hd__and4bb_2 _0957_ (.A_N(net115),
    .B_N(net221),
    .C(net116),
    .D(net117),
    .X(_0667_));
 sky130_fd_sc_hd__or3b_1 _0958_ (.A(_0648_),
    .B(_0654_),
    .C_N(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__a21o_1 _0959_ (.A1(net116),
    .A2(net117),
    .B1(net221),
    .X(_0669_));
 sky130_fd_sc_hd__and4b_1 _0960_ (.A_N(_0660_),
    .B(_0663_),
    .C(_0668_),
    .D(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _0961_ (.A0(net221),
    .A1(_0670_),
    .S(_0658_),
    .X(_0366_));
 sky130_fd_sc_hd__or2_1 _0962_ (.A(net116),
    .B(net118),
    .X(_0671_));
 sky130_fd_sc_hd__and3_1 _0963_ (.A(_0659_),
    .B(_0663_),
    .C(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _0964_ (.A0(net116),
    .A1(_0672_),
    .S(_0658_),
    .X(_0365_));
 sky130_fd_sc_hd__nor2_1 _0965_ (.A(net118),
    .B(_0498_),
    .Y(_0673_));
 sky130_fd_sc_hd__mux2_1 _0966_ (.A0(net118),
    .A1(_0673_),
    .S(_0658_),
    .X(_0364_));
 sky130_fd_sc_hd__nor3_1 _0967_ (.A(\state[2] ),
    .B(net312),
    .C(\state[0] ),
    .Y(_0674_));
 sky130_fd_sc_hd__nand2_2 _0968_ (.A(net299),
    .B(net313),
    .Y(_0675_));
 sky130_fd_sc_hd__or3_1 _0969_ (.A(_0489_),
    .B(net308),
    .C(net118),
    .X(_0676_));
 sky130_fd_sc_hd__and2_2 _0970_ (.A(net299),
    .B(_0654_),
    .X(_0677_));
 sky130_fd_sc_hd__nand3b_4 _0971_ (.A_N(net221),
    .B(net215),
    .C(net110),
    .Y(_0678_));
 sky130_fd_sc_hd__a2bb2o_1 _0972_ (.A1_N(_0676_),
    .A2_N(_0678_),
    .B1(net310),
    .B2(net113),
    .X(_0363_));
 sky130_fd_sc_hd__or3b_2 _0973_ (.A(net115),
    .B(net117),
    .C_N(net297),
    .X(_0679_));
 sky130_fd_sc_hd__a2bb2o_1 _0974_ (.A1_N(_0678_),
    .A2_N(_0679_),
    .B1(net179),
    .B2(net114),
    .X(_0362_));
 sky130_fd_sc_hd__or3b_2 _0975_ (.A(net115),
    .B(net118),
    .C_N(net249),
    .X(_0680_));
 sky130_fd_sc_hd__a2bb2o_1 _0976_ (.A1_N(_0678_),
    .A2_N(_0680_),
    .B1(net201),
    .B2(net111),
    .X(_0361_));
 sky130_fd_sc_hd__or3b_2 _0977_ (.A(net115),
    .B(net118),
    .C_N(net263),
    .X(_0681_));
 sky130_fd_sc_hd__a2bb2o_1 _0978_ (.A1_N(_0678_),
    .A2_N(_0681_),
    .B1(net173),
    .B2(net111),
    .X(_0360_));
 sky130_fd_sc_hd__or3b_2 _0979_ (.A(net115),
    .B(net118),
    .C_N(net219),
    .X(_0682_));
 sky130_fd_sc_hd__a2bb2o_1 _0980_ (.A1_N(_0678_),
    .A2_N(_0682_),
    .B1(net157),
    .B2(net111),
    .X(_0359_));
 sky130_fd_sc_hd__or3b_1 _0981_ (.A(net308),
    .B(net117),
    .C_N(net390),
    .X(_0683_));
 sky130_fd_sc_hd__a2bb2o_1 _0982_ (.A1_N(_0678_),
    .A2_N(_0683_),
    .B1(net347),
    .B2(net113),
    .X(_0358_));
 sky130_fd_sc_hd__or3b_1 _0983_ (.A(net115),
    .B(net118),
    .C_N(net256),
    .X(_0684_));
 sky130_fd_sc_hd__a2bb2o_1 _0984_ (.A1_N(_0678_),
    .A2_N(_0684_),
    .B1(net360),
    .B2(net112),
    .X(_0357_));
 sky130_fd_sc_hd__or3b_1 _0985_ (.A(net115),
    .B(net117),
    .C_N(net252),
    .X(_0685_));
 sky130_fd_sc_hd__a2bb2o_1 _0986_ (.A1_N(_0678_),
    .A2_N(net253),
    .B1(net145),
    .B2(net114),
    .X(_0356_));
 sky130_fd_sc_hd__nor2_1 _0987_ (.A(\byte_count[2] ),
    .B(net215),
    .Y(_0686_));
 sky130_fd_sc_hd__or2_4 _0988_ (.A(net221),
    .B(net215),
    .X(_0687_));
 sky130_fd_sc_hd__and3b_1 _0989_ (.A_N(net115),
    .B(net118),
    .C(net278),
    .X(_0688_));
 sky130_fd_sc_hd__and2_1 _0990_ (.A(net216),
    .B(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__a22o_1 _0991_ (.A1(net282),
    .A2(net111),
    .B1(net110),
    .B2(_0689_),
    .X(_0355_));
 sky130_fd_sc_hd__and3b_1 _0992_ (.A_N(net115),
    .B(net118),
    .C(net297),
    .X(_0690_));
 sky130_fd_sc_hd__and2_1 _0993_ (.A(net216),
    .B(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__a22o_1 _0994_ (.A1(net211),
    .A2(net111),
    .B1(net110),
    .B2(net217),
    .X(_0354_));
 sky130_fd_sc_hd__and3b_1 _0995_ (.A_N(net308),
    .B(net117),
    .C(net249),
    .X(_0692_));
 sky130_fd_sc_hd__and2_1 _0996_ (.A(net216),
    .B(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__a22o_1 _0997_ (.A1(net187),
    .A2(net113),
    .B1(net110),
    .B2(_0693_),
    .X(_0353_));
 sky130_fd_sc_hd__and3b_1 _0998_ (.A_N(net115),
    .B(net118),
    .C(net263),
    .X(_0694_));
 sky130_fd_sc_hd__and2_1 _0999_ (.A(net216),
    .B(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__a22o_1 _1000_ (.A1(net355),
    .A2(net112),
    .B1(net110),
    .B2(_0695_),
    .X(_0352_));
 sky130_fd_sc_hd__and3b_1 _1001_ (.A_N(net115),
    .B(net117),
    .C(net219),
    .X(_0696_));
 sky130_fd_sc_hd__and2_1 _1002_ (.A(net216),
    .B(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__a22o_1 _1003_ (.A1(net141),
    .A2(net113),
    .B1(net110),
    .B2(_0697_),
    .X(_0351_));
 sky130_fd_sc_hd__and3b_1 _1004_ (.A_N(net308),
    .B(net117),
    .C(net390),
    .X(_0698_));
 sky130_fd_sc_hd__and2_1 _1005_ (.A(net216),
    .B(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__a22o_1 _1006_ (.A1(net291),
    .A2(net114),
    .B1(net110),
    .B2(_0699_),
    .X(_0350_));
 sky130_fd_sc_hd__and3b_1 _1007_ (.A_N(\byte_count[3] ),
    .B(net118),
    .C(net256),
    .X(_0700_));
 sky130_fd_sc_hd__and2_1 _1008_ (.A(net216),
    .B(net257),
    .X(_0701_));
 sky130_fd_sc_hd__a22o_1 _1009_ (.A1(net225),
    .A2(net111),
    .B1(net110),
    .B2(_0701_),
    .X(_0349_));
 sky130_fd_sc_hd__and3b_1 _1010_ (.A_N(net115),
    .B(net229),
    .C(net252),
    .X(_0702_));
 sky130_fd_sc_hd__and2_1 _1011_ (.A(net216),
    .B(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__a22o_1 _1012_ (.A1(net306),
    .A2(net114),
    .B1(net110),
    .B2(_0703_),
    .X(_0348_));
 sky130_fd_sc_hd__nor2_1 _1013_ (.A(_0676_),
    .B(_0687_),
    .Y(_0704_));
 sky130_fd_sc_hd__a22o_1 _1014_ (.A1(net394),
    .A2(net113),
    .B1(_0677_),
    .B2(_0704_),
    .X(_0347_));
 sky130_fd_sc_hd__nor2_1 _1015_ (.A(_0679_),
    .B(_0687_),
    .Y(_0705_));
 sky130_fd_sc_hd__a22o_1 _1016_ (.A1(net245),
    .A2(net113),
    .B1(_0677_),
    .B2(_0705_),
    .X(_0346_));
 sky130_fd_sc_hd__nor2_1 _1017_ (.A(net250),
    .B(_0687_),
    .Y(_0706_));
 sky130_fd_sc_hd__a22o_1 _1018_ (.A1(net289),
    .A2(net114),
    .B1(net110),
    .B2(_0706_),
    .X(_0345_));
 sky130_fd_sc_hd__nor2_1 _1019_ (.A(net264),
    .B(_0687_),
    .Y(_0707_));
 sky130_fd_sc_hd__a22o_1 _1020_ (.A1(net366),
    .A2(net114),
    .B1(net110),
    .B2(_0707_),
    .X(_0344_));
 sky130_fd_sc_hd__nor2_1 _1021_ (.A(_0682_),
    .B(_0687_),
    .Y(_0708_));
 sky130_fd_sc_hd__a22o_1 _1022_ (.A1(net365),
    .A2(net111),
    .B1(net110),
    .B2(_0708_),
    .X(_0343_));
 sky130_fd_sc_hd__nor2_2 _1023_ (.A(_0683_),
    .B(_0687_),
    .Y(_0434_));
 sky130_fd_sc_hd__a22o_1 _1024_ (.A1(net199),
    .A2(net112),
    .B1(net110),
    .B2(_0434_),
    .X(_0342_));
 sky130_fd_sc_hd__nor2_1 _1025_ (.A(_0684_),
    .B(_0687_),
    .Y(_0435_));
 sky130_fd_sc_hd__a22o_1 _1026_ (.A1(net284),
    .A2(net112),
    .B1(net110),
    .B2(_0435_),
    .X(_0341_));
 sky130_fd_sc_hd__nor2_2 _1027_ (.A(_0685_),
    .B(_0687_),
    .Y(_0436_));
 sky130_fd_sc_hd__a22o_1 _1028_ (.A1(net247),
    .A2(net113),
    .B1(net110),
    .B2(_0436_),
    .X(_0340_));
 sky130_fd_sc_hd__and2_2 _1029_ (.A(net299),
    .B(_0661_),
    .X(_0437_));
 sky130_fd_sc_hd__and3b_4 _1030_ (.A_N(net221),
    .B(net116),
    .C(net109),
    .X(_0438_));
 sky130_fd_sc_hd__nand3b_4 _1031_ (.A_N(net221),
    .B(net116),
    .C(net109),
    .Y(_0439_));
 sky130_fd_sc_hd__a22o_1 _1032_ (.A1(net369),
    .A2(net111),
    .B1(net279),
    .B2(_0438_),
    .X(_0339_));
 sky130_fd_sc_hd__a22o_1 _1033_ (.A1(net371),
    .A2(net111),
    .B1(_0690_),
    .B2(_0438_),
    .X(_0338_));
 sky130_fd_sc_hd__a22o_1 _1034_ (.A1(net388),
    .A2(net113),
    .B1(_0692_),
    .B2(_0438_),
    .X(_0337_));
 sky130_fd_sc_hd__a22o_1 _1035_ (.A1(net233),
    .A2(net112),
    .B1(_0694_),
    .B2(_0438_),
    .X(_0336_));
 sky130_fd_sc_hd__a22o_1 _1036_ (.A1(net193),
    .A2(net113),
    .B1(_0696_),
    .B2(_0438_),
    .X(_0335_));
 sky130_fd_sc_hd__a22o_1 _1037_ (.A1(net207),
    .A2(net113),
    .B1(_0698_),
    .B2(_0438_),
    .X(_0334_));
 sky130_fd_sc_hd__a22o_1 _1038_ (.A1(net161),
    .A2(net112),
    .B1(net257),
    .B2(_0438_),
    .X(_0333_));
 sky130_fd_sc_hd__a22o_1 _1039_ (.A1(net398),
    .A2(net113),
    .B1(_0702_),
    .B2(_0438_),
    .X(_0332_));
 sky130_fd_sc_hd__a2bb2o_1 _1040_ (.A1_N(_0676_),
    .A2_N(_0439_),
    .B1(net374),
    .B2(net113),
    .X(_0331_));
 sky130_fd_sc_hd__a2bb2o_1 _1041_ (.A1_N(_0679_),
    .A2_N(_0439_),
    .B1(net205),
    .B2(net114),
    .X(_0330_));
 sky130_fd_sc_hd__a2bb2o_1 _1042_ (.A1_N(_0680_),
    .A2_N(_0439_),
    .B1(net177),
    .B2(net114),
    .X(_0329_));
 sky130_fd_sc_hd__a2bb2o_1 _1043_ (.A1_N(net264),
    .A2_N(_0439_),
    .B1(net185),
    .B2(net114),
    .X(_0328_));
 sky130_fd_sc_hd__a2bb2o_1 _1044_ (.A1_N(_0682_),
    .A2_N(_0439_),
    .B1(net163),
    .B2(net112),
    .X(_0327_));
 sky130_fd_sc_hd__a2bb2o_1 _1045_ (.A1_N(_0683_),
    .A2_N(_0439_),
    .B1(net367),
    .B2(net113),
    .X(_0326_));
 sky130_fd_sc_hd__a2bb2o_1 _1046_ (.A1_N(_0684_),
    .A2_N(_0439_),
    .B1(net153),
    .B2(net112),
    .X(_0325_));
 sky130_fd_sc_hd__a2bb2o_1 _1047_ (.A1_N(net253),
    .A2_N(_0439_),
    .B1(net351),
    .B2(net114),
    .X(_0324_));
 sky130_fd_sc_hd__a22o_1 _1048_ (.A1(net235),
    .A2(net111),
    .B1(_0689_),
    .B2(net109),
    .X(_0323_));
 sky130_fd_sc_hd__a22o_1 _1049_ (.A1(net337),
    .A2(net111),
    .B1(net217),
    .B2(net109),
    .X(_0322_));
 sky130_fd_sc_hd__a22o_1 _1050_ (.A1(net181),
    .A2(net114),
    .B1(_0693_),
    .B2(net109),
    .X(_0321_));
 sky130_fd_sc_hd__a22o_1 _1051_ (.A1(net169),
    .A2(net111),
    .B1(_0695_),
    .B2(net109),
    .X(_0320_));
 sky130_fd_sc_hd__a22o_1 _1052_ (.A1(net400),
    .A2(net112),
    .B1(_0697_),
    .B2(net109),
    .X(_0319_));
 sky130_fd_sc_hd__a22o_1 _1053_ (.A1(net261),
    .A2(net113),
    .B1(_0699_),
    .B2(net109),
    .X(_0318_));
 sky130_fd_sc_hd__a22o_1 _1054_ (.A1(net421),
    .A2(net111),
    .B1(_0701_),
    .B2(net109),
    .X(_0317_));
 sky130_fd_sc_hd__a22o_1 _1055_ (.A1(net266),
    .A2(net114),
    .B1(_0703_),
    .B2(net109),
    .X(_0316_));
 sky130_fd_sc_hd__a22o_1 _1056_ (.A1(net335),
    .A2(net114),
    .B1(_0704_),
    .B2(net109),
    .X(_0315_));
 sky130_fd_sc_hd__a22o_1 _1057_ (.A1(net171),
    .A2(net114),
    .B1(_0705_),
    .B2(net109),
    .X(_0314_));
 sky130_fd_sc_hd__a22o_1 _1058_ (.A1(net293),
    .A2(net113),
    .B1(_0706_),
    .B2(_0437_),
    .X(_0313_));
 sky130_fd_sc_hd__a22o_1 _1059_ (.A1(net330),
    .A2(net114),
    .B1(_0707_),
    .B2(net300),
    .X(_0312_));
 sky130_fd_sc_hd__a22o_1 _1060_ (.A1(net223),
    .A2(net111),
    .B1(_0708_),
    .B2(net109),
    .X(_0311_));
 sky130_fd_sc_hd__a22o_1 _1061_ (.A1(net203),
    .A2(net113),
    .B1(_0434_),
    .B2(net300),
    .X(_0310_));
 sky130_fd_sc_hd__a22o_1 _1062_ (.A1(net227),
    .A2(_0675_),
    .B1(_0435_),
    .B2(net109),
    .X(_0309_));
 sky130_fd_sc_hd__a22o_1 _1063_ (.A1(net209),
    .A2(net111),
    .B1(_0436_),
    .B2(net109),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _1064_ (.A0(net278),
    .A1(net373),
    .S(net112),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _1065_ (.A0(net297),
    .A1(net387),
    .S(net112),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _1066_ (.A0(net249),
    .A1(net379),
    .S(net112),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _1067_ (.A0(net263),
    .A1(net358),
    .S(net112),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _1068_ (.A0(net219),
    .A1(net393),
    .S(_0675_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _1069_ (.A0(net506),
    .A1(net377),
    .S(net111),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _1070_ (.A0(net256),
    .A1(net384),
    .S(net112),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _1071_ (.A0(net252),
    .A1(net364),
    .S(net112),
    .X(_0300_));
 sky130_fd_sc_hd__and2b_1 _1072_ (.A_N(net299),
    .B(net313),
    .X(_0440_));
 sky130_fd_sc_hd__nor2_1 _1073_ (.A(_0648_),
    .B(net313),
    .Y(_0441_));
 sky130_fd_sc_hd__a211o_1 _1074_ (.A1(_0648_),
    .A2(net242),
    .B1(_0440_),
    .C1(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__nor3b_4 _1075_ (.A(net115),
    .B(net221),
    .C_N(_0648_),
    .Y(_0443_));
 sky130_fd_sc_hd__mux4_1 _1076_ (.A0(net34),
    .A1(net11),
    .A2(net20),
    .A3(net29),
    .S0(net117),
    .S1(net116),
    .X(_0444_));
 sky130_fd_sc_hd__and2_1 _1077_ (.A(_0443_),
    .B(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _1078_ (.A0(_0445_),
    .A1(net149),
    .S(net243),
    .X(_0299_));
 sky130_fd_sc_hd__mux4_1 _1079_ (.A0(net33),
    .A1(net10),
    .A2(net19),
    .A3(net28),
    .S0(net117),
    .S1(net116),
    .X(_0446_));
 sky130_fd_sc_hd__and2_1 _1080_ (.A(_0443_),
    .B(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _1081_ (.A0(_0447_),
    .A1(net155),
    .S(net243),
    .X(_0298_));
 sky130_fd_sc_hd__mux4_1 _1082_ (.A0(net32),
    .A1(net9),
    .A2(net18),
    .A3(net26),
    .S0(net117),
    .S1(net116),
    .X(_0448_));
 sky130_fd_sc_hd__and2_1 _1083_ (.A(_0443_),
    .B(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _1084_ (.A0(_0449_),
    .A1(net239),
    .S(_0442_),
    .X(_0297_));
 sky130_fd_sc_hd__mux4_1 _1085_ (.A0(net31),
    .A1(net8),
    .A2(net17),
    .A3(net25),
    .S0(net117),
    .S1(net116),
    .X(_0450_));
 sky130_fd_sc_hd__and2_1 _1086_ (.A(_0443_),
    .B(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _1087_ (.A0(_0451_),
    .A1(net276),
    .S(net243),
    .X(_0296_));
 sky130_fd_sc_hd__mux4_1 _1088_ (.A0(net30),
    .A1(net7),
    .A2(net15),
    .A3(net24),
    .S0(net117),
    .S1(net116),
    .X(_0452_));
 sky130_fd_sc_hd__and2_1 _1089_ (.A(_0443_),
    .B(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _1090_ (.A0(_0453_),
    .A1(net349),
    .S(net243),
    .X(_0295_));
 sky130_fd_sc_hd__mux4_1 _1091_ (.A0(net27),
    .A1(net6),
    .A2(net14),
    .A3(net23),
    .S0(net118),
    .S1(net116),
    .X(_0454_));
 sky130_fd_sc_hd__and2_1 _1092_ (.A(_0443_),
    .B(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _1093_ (.A0(_0455_),
    .A1(net270),
    .S(net243),
    .X(_0294_));
 sky130_fd_sc_hd__mux4_1 _1094_ (.A0(net16),
    .A1(net36),
    .A2(net13),
    .A3(net22),
    .S0(net117),
    .S1(net116),
    .X(_0456_));
 sky130_fd_sc_hd__and2_1 _1095_ (.A(_0443_),
    .B(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _1096_ (.A0(_0457_),
    .A1(net195),
    .S(_0442_),
    .X(_0293_));
 sky130_fd_sc_hd__mux4_1 _1097_ (.A0(net5),
    .A1(net35),
    .A2(net12),
    .A3(net21),
    .S0(net118),
    .S1(net116),
    .X(_0458_));
 sky130_fd_sc_hd__and2_1 _1098_ (.A(_0443_),
    .B(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _1099_ (.A0(_0459_),
    .A1(net143),
    .S(net243),
    .X(_0292_));
 sky130_fd_sc_hd__or4b_1 _1100_ (.A(net115),
    .B(net116),
    .C(net117),
    .D_N(net221),
    .X(_0460_));
 sky130_fd_sc_hd__and4b_1 _1101_ (.A_N(net391),
    .B(net241),
    .C(_0648_),
    .D(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__a21o_1 _1102_ (.A1(net391),
    .A2(_0441_),
    .B1(_0461_),
    .X(_0291_));
 sky130_fd_sc_hd__nand2_4 _1103_ (.A(_0667_),
    .B(net110),
    .Y(_0462_));
 sky130_fd_sc_hd__mux2_1 _1104_ (.A0(net278),
    .A1(net404),
    .S(net108),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _1105_ (.A0(net297),
    .A1(net460),
    .S(net107),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _1106_ (.A0(net249),
    .A1(net468),
    .S(net107),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _1107_ (.A0(net263),
    .A1(net462),
    .S(net107),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _1108_ (.A0(net219),
    .A1(net461),
    .S(net108),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _1109_ (.A0(net390),
    .A1(net440),
    .S(net107),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _1110_ (.A0(net256),
    .A1(net423),
    .S(net108),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _1111_ (.A0(net252),
    .A1(net441),
    .S(net107),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _1112_ (.A0(net310),
    .A1(net86),
    .S(net108),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _1113_ (.A0(net179),
    .A1(net85),
    .S(net108),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _1114_ (.A0(net201),
    .A1(net84),
    .S(net107),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _1115_ (.A0(net173),
    .A1(net83),
    .S(net107),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _1116_ (.A0(net157),
    .A1(net81),
    .S(net107),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _1117_ (.A0(net347),
    .A1(net80),
    .S(net108),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _1118_ (.A0(net360),
    .A1(net79),
    .S(net108),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _1119_ (.A0(net145),
    .A1(net78),
    .S(net107),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _1120_ (.A0(net282),
    .A1(net323),
    .S(net107),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _1121_ (.A0(net211),
    .A1(net76),
    .S(net107),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _1122_ (.A0(net187),
    .A1(net75),
    .S(net108),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _1123_ (.A0(net355),
    .A1(net359),
    .S(net107),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _1124_ (.A0(net141),
    .A1(net73),
    .S(net108),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _1125_ (.A0(net291),
    .A1(net321),
    .S(net107),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _1126_ (.A0(net225),
    .A1(net231),
    .S(net107),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _1127_ (.A0(net306),
    .A1(net101),
    .S(net107),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _1128_ (.A0(net394),
    .A1(net100),
    .S(_0462_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _1129_ (.A0(net245),
    .A1(net339),
    .S(_0462_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _1130_ (.A0(net289),
    .A1(net302),
    .S(net108),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _1131_ (.A0(net366),
    .A1(net376),
    .S(net108),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _1132_ (.A0(net365),
    .A1(net372),
    .S(net108),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _1133_ (.A0(net199),
    .A1(net304),
    .S(net107),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _1134_ (.A0(net284),
    .A1(net316),
    .S(net108),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _1135_ (.A0(net247),
    .A1(net268),
    .S(net108),
    .X(_0259_));
 sky130_fd_sc_hd__and4b_1 _1136_ (.A_N(net373),
    .B(net387),
    .C(net379),
    .D(net358),
    .X(_0463_));
 sky130_fd_sc_hd__and4b_1 _1137_ (.A_N(net393),
    .B(net377),
    .C(net384),
    .D(net364),
    .X(_0464_));
 sky130_fd_sc_hd__nand2_1 _1138_ (.A(_0463_),
    .B(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__a21oi_1 _1139_ (.A1(_0463_),
    .A2(_0464_),
    .B1(_0662_),
    .Y(_0466_));
 sky130_fd_sc_hd__nand2_1 _1140_ (.A(net299),
    .B(_0667_),
    .Y(_0467_));
 sky130_fd_sc_hd__or4_4 _1141_ (.A(net411),
    .B(_0498_),
    .C(_0466_),
    .D(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _1142_ (.A0(net369),
    .A1(net62),
    .S(net106),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _1143_ (.A0(net371),
    .A1(net385),
    .S(net106),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _1144_ (.A0(net388),
    .A1(net59),
    .S(net105),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _1145_ (.A0(net233),
    .A1(net58),
    .S(net106),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _1146_ (.A0(net193),
    .A1(net213),
    .S(net105),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _1147_ (.A0(net207),
    .A1(net56),
    .S(net106),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _1148_ (.A0(net161),
    .A1(net55),
    .S(net106),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _1149_ (.A0(net398),
    .A1(net54),
    .S(net105),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _1150_ (.A0(net374),
    .A1(net53),
    .S(net105),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _1151_ (.A0(net205),
    .A1(net52),
    .S(net105),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _1152_ (.A0(net177),
    .A1(net51),
    .S(net105),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _1153_ (.A0(net185),
    .A1(net50),
    .S(net105),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _1154_ (.A0(net163),
    .A1(net48),
    .S(net106),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _1155_ (.A0(net367),
    .A1(net47),
    .S(net105),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _1156_ (.A0(net153),
    .A1(net46),
    .S(net106),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _1157_ (.A0(net351),
    .A1(net45),
    .S(net105),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _1158_ (.A0(net235),
    .A1(net44),
    .S(net106),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _1159_ (.A0(net337),
    .A1(net43),
    .S(net106),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _1160_ (.A0(net181),
    .A1(net42),
    .S(net105),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _1161_ (.A0(net169),
    .A1(net41),
    .S(net106),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _1162_ (.A0(net400),
    .A1(net40),
    .S(net106),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _1163_ (.A0(net261),
    .A1(net328),
    .S(net105),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _1164_ (.A0(net421),
    .A1(net69),
    .S(net105),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _1165_ (.A0(net266),
    .A1(net295),
    .S(net105),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _1166_ (.A0(net335),
    .A1(net353),
    .S(net105),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _1167_ (.A0(net171),
    .A1(net66),
    .S(net105),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _1168_ (.A0(net293),
    .A1(net319),
    .S(net105),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _1169_ (.A0(net330),
    .A1(net341),
    .S(_0468_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _1170_ (.A0(net223),
    .A1(net63),
    .S(net106),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _1171_ (.A0(net203),
    .A1(net60),
    .S(_0468_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _1172_ (.A0(net227),
    .A1(net286),
    .S(net106),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _1173_ (.A0(net209),
    .A1(net237),
    .S(net106),
    .X(_0227_));
 sky130_fd_sc_hd__a211oi_1 _1174_ (.A1(net299),
    .A2(_0667_),
    .B1(net411),
    .C1(_0498_),
    .Y(_0469_));
 sky130_fd_sc_hd__o22a_1 _1175_ (.A1(_0499_),
    .A2(_0650_),
    .B1(_0652_),
    .B2(\state[2] ),
    .X(_0470_));
 sky130_fd_sc_hd__a311o_1 _1176_ (.A1(net299),
    .A2(_0667_),
    .A3(_0466_),
    .B1(_0469_),
    .C1(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__a21bo_1 _1177_ (.A1(net407),
    .A2(_0471_),
    .B1_N(net108),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _1178_ (.A0(net109),
    .A1(_0466_),
    .S(_0667_),
    .X(_0472_));
 sky130_fd_sc_hd__or3_2 _1179_ (.A(_0651_),
    .B(_0461_),
    .C(_0469_),
    .X(_0473_));
 sky130_fd_sc_hd__or3_1 _1180_ (.A(net418),
    .B(_0472_),
    .C(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__a21bo_1 _1181_ (.A1(net471),
    .A2(_0474_),
    .B1_N(net106),
    .X(_0225_));
 sky130_fd_sc_hd__a32o_1 _1182_ (.A1(net356),
    .A2(_0544_),
    .A3(net414),
    .B1(_0567_),
    .B2(net241),
    .X(_0224_));
 sky130_fd_sc_hd__nor2_1 _1183_ (.A(_0440_),
    .B(_0473_),
    .Y(_0475_));
 sky130_fd_sc_hd__nor2_1 _1184_ (.A(_0662_),
    .B(_0465_),
    .Y(_0476_));
 sky130_fd_sc_hd__or3_1 _1185_ (.A(_0653_),
    .B(_0654_),
    .C(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__a211o_1 _1186_ (.A1(_0475_),
    .A2(_0477_),
    .B1(_0651_),
    .C1(_0461_),
    .X(_0223_));
 sky130_fd_sc_hd__and4bb_1 _1187_ (.A_N(net377),
    .B_N(net364),
    .C(net384),
    .D(net393),
    .X(_0478_));
 sky130_fd_sc_hd__and4bb_1 _1188_ (.A_N(net387),
    .B_N(net358),
    .C(net379),
    .D(net373),
    .X(_0479_));
 sky130_fd_sc_hd__a31o_1 _1189_ (.A1(net412),
    .A2(_0478_),
    .A3(_0479_),
    .B1(_0653_),
    .X(_0480_));
 sky130_fd_sc_hd__or4b_1 _1190_ (.A(net263),
    .B(net390),
    .C(net252),
    .D_N(\uart_rx_inst.o_data[3] ),
    .X(_0481_));
 sky130_fd_sc_hd__nor3_1 _1191_ (.A(_0489_),
    .B(net297),
    .C(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__and4b_1 _1192_ (.A_N(\uart_rx_inst.o_data[3] ),
    .B(net390),
    .C(net252),
    .D(net263),
    .X(_0483_));
 sky130_fd_sc_hd__a31o_1 _1193_ (.A1(_0489_),
    .A2(net297),
    .A3(_0483_),
    .B1(_0482_),
    .X(_0484_));
 sky130_fd_sc_hd__a41o_1 _1194_ (.A1(net249),
    .A2(net256),
    .A3(net313),
    .A4(_0484_),
    .B1(_0480_),
    .X(_0485_));
 sky130_fd_sc_hd__a22o_1 _1195_ (.A1(net312),
    .A2(_0473_),
    .B1(_0475_),
    .B2(_0485_),
    .X(_0222_));
 sky130_fd_sc_hd__a21bo_1 _1196_ (.A1(_0478_),
    .A2(_0479_),
    .B1_N(_0465_),
    .X(_0486_));
 sky130_fd_sc_hd__a32o_1 _1197_ (.A1(net412),
    .A2(_0475_),
    .A3(_0486_),
    .B1(_0473_),
    .B2(net418),
    .X(_0221_));
 sky130_fd_sc_hd__nand2b_1 _1198_ (.A_N(net165),
    .B(net1),
    .Y(_0487_));
 sky130_fd_sc_hd__a21oi_1 _1199_ (.A1(_0500_),
    .A2(_0487_),
    .B1(net333),
    .Y(_0001_));
 sky130_fd_sc_hd__a31oi_1 _1200_ (.A1(net356),
    .A2(_0544_),
    .A3(_0600_),
    .B1(_0546_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _1201_ (.A(net127),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _1202_ (.A(net127),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _1203_ (.A(net128),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _1204_ (.A(net122),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _1205_ (.A(net128),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _1206_ (.A(net119),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _1207_ (.A(net123),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _1208_ (.A(net133),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _1209_ (.A(net119),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _1210_ (.A(net133),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1211_ (.A(net133),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _1212_ (.A(net129),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _1213_ (.A(net129),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _1214_ (.A(net130),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _1215_ (.A(net129),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _1216_ (.A(net132),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _1217_ (.A(net123),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _1218_ (.A(net120),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _1219_ (.A(net133),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _1220_ (.A(net123),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _1221_ (.A(net120),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1222_ (.A(net129),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _1223_ (.A(net120),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1224_ (.A(net130),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1225_ (.A(net123),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1226_ (.A(net133),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _1227_ (.A(net129),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _1228_ (.A(net129),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _1229_ (.A(net133),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _1230_ (.A(net133),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1231_ (.A(net124),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _1232_ (.A(net123),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1233_ (.A(net131),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _1234_ (.A(net121),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _1235_ (.A(net133),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _1236_ (.A(net119),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1237_ (.A(net119),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _1238_ (.A(net131),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _1239_ (.A(net124),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _1240_ (.A(net121),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _1241_ (.A(net121),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _1242_ (.A(net133),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _1243_ (.A(net133),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _1244_ (.A(net132),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _1245_ (.A(net124),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _1246_ (.A(net127),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _1247_ (.A(net120),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _1248_ (.A(net129),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _1249_ (.A(net131),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _1250_ (.A(net121),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _1251_ (.A(net132),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _1252_ (.A(net120),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _1253_ (.A(net119),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _1254_ (.A(net127),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _1255_ (.A(net124),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _1256_ (.A(net125),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _1257_ (.A(net119),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _1258_ (.A(net119),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _1259_ (.A(net119),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _1260_ (.A(net132),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _1261_ (.A(net132),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _1262_ (.A(net121),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _1263_ (.A(net132),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _1264_ (.A(net127),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _1265_ (.A(net124),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _1266_ (.A(net120),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _1267_ (.A(net119),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _1268_ (.A(net121),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _1269_ (.A(net131),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _1270_ (.A(net128),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _1271_ (.A(net128),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _1272_ (.A(net128),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _1273_ (.A(net128),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _1274_ (.A(net129),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _1275_ (.A(net127),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _1276_ (.A(net127),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _1277_ (.A(net127),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _1278_ (.A(net129),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _1279_ (.A(net125),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _1280_ (.A(net125),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _1281_ (.A(net122),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _1282_ (.A(net122),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _1283_ (.A(net122),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _1284_ (.A(net121),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _1285_ (.A(net122),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _1286_ (.A(net122),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _1287_ (.A(net119),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _1288_ (.A(net123),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _1289_ (.A(net134),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _1290_ (.A(net119),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _1291_ (.A(net134),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _1292_ (.A(net134),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _1293_ (.A(net129),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _1294_ (.A(net127),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _1295_ (.A(net130),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _1296_ (.A(net120),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _1297_ (.A(net132),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _1298_ (.A(net125),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _1299_ (.A(net119),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _1300_ (.A(net132),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _1301_ (.A(net120),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _1302_ (.A(net120),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _1303_ (.A(net127),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _1304_ (.A(net123),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _1305_ (.A(net131),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _1306_ (.A(net123),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _1307_ (.A(net134),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _1308_ (.A(net129),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _1309_ (.A(net129),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _1310_ (.A(net131),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _1311_ (.A(net131),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _1312_ (.A(net123),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _1313_ (.A(net131),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _1314_ (.A(net131),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _1315_ (.A(net121),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _1316_ (.A(net132),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _1317_ (.A(net120),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _1318_ (.A(net119),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _1319_ (.A(net131),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _1320_ (.A(net124),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _1321_ (.A(net121),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _1322_ (.A(net121),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _1323_ (.A(net134),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _1324_ (.A(net134),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _1325_ (.A(net132),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _1326_ (.A(net132),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _1327_ (.A(net127),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _1328_ (.A(net120),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _1329_ (.A(net129),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _1330_ (.A(net131),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _1331_ (.A(net121),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _1332_ (.A(net132),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _1333_ (.A(net120),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _1334_ (.A(net119),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _1335_ (.A(net127),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _1336_ (.A(net123),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _1337_ (.A(net125),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _1338_ (.A(net119),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _1339_ (.A(net119),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _1340_ (.A(net135),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _1341_ (.A(net131),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _1342_ (.A(net131),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _1343_ (.A(net121),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _1344_ (.A(net121),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _1345_ (.A(net127),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _1346_ (.A(net121),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _1347_ (.A(net129),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _1348_ (.A(net125),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _1349_ (.A(net124),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _1350_ (.A(net124),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _1351_ (.A(net124),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _1352_ (.A(net124),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _1353_ (.A(net125),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _1354_ (.A(net125),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _1355_ (.A(net125),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _1356_ (.A(net126),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _1357_ (.A(net126),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _1358_ (.A(net126),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _1359_ (.A(net126),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _1360_ (.A(net126),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _1361_ (.A(net124),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _1362_ (.A(net126),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _1363_ (.A(net124),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _1364_ (.A(net126),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _1365_ (.A(net123),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _1366_ (.A(net123),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _1367_ (.A(net123),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _1368_ (.A(net123),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _1369_ (.A(net125),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _1370_ (.A(net125),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _1371_ (.A(net125),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _1372_ (.A(net125),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _1373_ (.A(net122),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _1374_ (.A(net120),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _1375_ (.A(net120),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _1376_ (.A(net123),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _1377_ (.A(net122),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _1378_ (.A(net128),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _1379_ (.A(net128),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _1380_ (.A(net128),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _1381_ (.A(net129),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _1382_ (.A(net127),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _1383_ (.A(net127),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _1384_ (.A(net127),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _1385_ (.A(net129),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _1386_ (.A(net130),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _1387_ (.A(net121),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _1388_ (.A(net130),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _1389_ (.A(net128),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _1390_ (.A(net133),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _1391_ (.A(net131),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _1392_ (.A(net131),
    .Y(_0195_));
 sky130_fd_sc_hd__inv_2 _1393_ (.A(net133),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_2 _1394_ (.A(net133),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_2 _1395_ (.A(net133),
    .Y(_0198_));
 sky130_fd_sc_hd__inv_2 _1396_ (.A(net133),
    .Y(_0199_));
 sky130_fd_sc_hd__inv_2 _1397_ (.A(net133),
    .Y(_0200_));
 sky130_fd_sc_hd__inv_2 _1398_ (.A(net130),
    .Y(_0201_));
 sky130_fd_sc_hd__inv_2 _1399_ (.A(net130),
    .Y(_0202_));
 sky130_fd_sc_hd__inv_2 _1400_ (.A(net130),
    .Y(_0203_));
 sky130_fd_sc_hd__inv_2 _1401_ (.A(net130),
    .Y(_0204_));
 sky130_fd_sc_hd__inv_2 _1402_ (.A(net128),
    .Y(_0205_));
 sky130_fd_sc_hd__inv_2 _1403_ (.A(net130),
    .Y(_0206_));
 sky130_fd_sc_hd__inv_2 _1404_ (.A(net131),
    .Y(_0207_));
 sky130_fd_sc_hd__inv_2 _1405_ (.A(net132),
    .Y(_0208_));
 sky130_fd_sc_hd__inv_2 _1406_ (.A(net130),
    .Y(_0209_));
 sky130_fd_sc_hd__inv_2 _1407_ (.A(net130),
    .Y(_0210_));
 sky130_fd_sc_hd__inv_2 _1408_ (.A(net130),
    .Y(_0211_));
 sky130_fd_sc_hd__inv_2 _1409_ (.A(net130),
    .Y(_0212_));
 sky130_fd_sc_hd__inv_2 _1410_ (.A(net122),
    .Y(_0213_));
 sky130_fd_sc_hd__inv_2 _1411_ (.A(net125),
    .Y(_0214_));
 sky130_fd_sc_hd__inv_2 _1412_ (.A(net125),
    .Y(_0215_));
 sky130_fd_sc_hd__inv_2 _1413_ (.A(net125),
    .Y(_0216_));
 sky130_fd_sc_hd__inv_2 _1414_ (.A(net120),
    .Y(_0217_));
 sky130_fd_sc_hd__inv_2 _1415_ (.A(net120),
    .Y(_0218_));
 sky130_fd_sc_hd__inv_2 _1416_ (.A(net135),
    .Y(_0219_));
 sky130_fd_sc_hd__inv_2 _1417_ (.A(net123),
    .Y(_0220_));
 sky130_fd_sc_hd__dfrtp_1 _1418_ (.CLK(clknet_leaf_2_clk),
    .D(_0221_),
    .RESET_B(_0003_),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1419_ (.CLK(clknet_leaf_23_clk),
    .D(_0222_),
    .RESET_B(_0004_),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1420_ (.CLK(clknet_leaf_22_clk),
    .D(_0223_),
    .RESET_B(_0005_),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfstp_1 _1421_ (.CLK(clknet_leaf_16_clk),
    .D(net415),
    .SET_B(_0006_),
    .Q(\uart_tx_inst.o_ready ));
 sky130_fd_sc_hd__dfrtp_4 _1422_ (.CLK(clknet_leaf_2_clk),
    .D(_0225_),
    .RESET_B(_0007_),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_2 _1423_ (.CLK(clknet_leaf_15_clk),
    .D(net408),
    .RESET_B(_0008_),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 _1424_ (.CLK(clknet_leaf_27_clk),
    .D(net238),
    .RESET_B(_0009_),
    .Q(net38));
 sky130_fd_sc_hd__dfrtp_1 _1425_ (.CLK(clknet_leaf_5_clk),
    .D(net287),
    .RESET_B(_0010_),
    .Q(net49));
 sky130_fd_sc_hd__dfrtp_2 _1426_ (.CLK(clknet_leaf_12_clk),
    .D(net204),
    .RESET_B(_0011_),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_1 _1427_ (.CLK(clknet_leaf_27_clk),
    .D(net224),
    .RESET_B(_0012_),
    .Q(net63));
 sky130_fd_sc_hd__dfrtp_1 _1428_ (.CLK(clknet_leaf_12_clk),
    .D(net342),
    .RESET_B(_0013_),
    .Q(net64));
 sky130_fd_sc_hd__dfrtp_1 _1429_ (.CLK(clknet_leaf_12_clk),
    .D(net320),
    .RESET_B(_0014_),
    .Q(net65));
 sky130_fd_sc_hd__dfrtp_1 _1430_ (.CLK(clknet_leaf_19_clk),
    .D(net172),
    .RESET_B(_0015_),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_1 _1431_ (.CLK(clknet_leaf_20_clk),
    .D(net354),
    .RESET_B(_0016_),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _1432_ (.CLK(clknet_leaf_17_clk),
    .D(net296),
    .RESET_B(_0017_),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_1 _1433_ (.CLK(clknet_leaf_18_clk),
    .D(net422),
    .RESET_B(_0018_),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _1434_ (.CLK(clknet_leaf_11_clk),
    .D(net329),
    .RESET_B(_0019_),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_1 _1435_ (.CLK(clknet_leaf_5_clk),
    .D(net401),
    .RESET_B(_0020_),
    .Q(net40));
 sky130_fd_sc_hd__dfrtp_1 _1436_ (.CLK(clknet_leaf_0_clk),
    .D(net170),
    .RESET_B(_0021_),
    .Q(net41));
 sky130_fd_sc_hd__dfrtp_1 _1437_ (.CLK(clknet_leaf_12_clk),
    .D(net182),
    .RESET_B(_0022_),
    .Q(net42));
 sky130_fd_sc_hd__dfrtp_1 _1438_ (.CLK(clknet_leaf_6_clk),
    .D(net338),
    .RESET_B(_0023_),
    .Q(net43));
 sky130_fd_sc_hd__dfrtp_1 _1439_ (.CLK(clknet_leaf_1_clk),
    .D(net236),
    .RESET_B(_0024_),
    .Q(net44));
 sky130_fd_sc_hd__dfrtp_1 _1440_ (.CLK(clknet_leaf_18_clk),
    .D(net352),
    .RESET_B(_0025_),
    .Q(net45));
 sky130_fd_sc_hd__dfrtp_1 _1441_ (.CLK(clknet_leaf_1_clk),
    .D(net154),
    .RESET_B(_0026_),
    .Q(net46));
 sky130_fd_sc_hd__dfrtp_1 _1442_ (.CLK(clknet_leaf_16_clk),
    .D(net368),
    .RESET_B(_0027_),
    .Q(net47));
 sky130_fd_sc_hd__dfrtp_1 _1443_ (.CLK(clknet_leaf_6_clk),
    .D(net164),
    .RESET_B(_0028_),
    .Q(net48));
 sky130_fd_sc_hd__dfrtp_1 _1444_ (.CLK(clknet_leaf_12_clk),
    .D(net186),
    .RESET_B(_0029_),
    .Q(net50));
 sky130_fd_sc_hd__dfrtp_1 _1445_ (.CLK(clknet_leaf_19_clk),
    .D(net178),
    .RESET_B(_0030_),
    .Q(net51));
 sky130_fd_sc_hd__dfrtp_1 _1446_ (.CLK(clknet_leaf_19_clk),
    .D(net206),
    .RESET_B(_0031_),
    .Q(net52));
 sky130_fd_sc_hd__dfrtp_1 _1447_ (.CLK(clknet_leaf_13_clk),
    .D(net375),
    .RESET_B(_0032_),
    .Q(net53));
 sky130_fd_sc_hd__dfrtp_1 _1448_ (.CLK(clknet_leaf_12_clk),
    .D(net399),
    .RESET_B(_0033_),
    .Q(net54));
 sky130_fd_sc_hd__dfrtp_1 _1449_ (.CLK(clknet_leaf_6_clk),
    .D(net162),
    .RESET_B(_0034_),
    .Q(net55));
 sky130_fd_sc_hd__dfrtp_1 _1450_ (.CLK(clknet_leaf_5_clk),
    .D(net208),
    .RESET_B(_0035_),
    .Q(net56));
 sky130_fd_sc_hd__dfrtp_2 _1451_ (.CLK(clknet_leaf_10_clk),
    .D(net214),
    .RESET_B(_0036_),
    .Q(net57));
 sky130_fd_sc_hd__dfrtp_1 _1452_ (.CLK(clknet_leaf_24_clk),
    .D(net234),
    .RESET_B(_0037_),
    .Q(net58));
 sky130_fd_sc_hd__dfrtp_1 _1453_ (.CLK(clknet_leaf_12_clk),
    .D(net389),
    .RESET_B(_0038_),
    .Q(net59));
 sky130_fd_sc_hd__dfrtp_1 _1454_ (.CLK(clknet_leaf_0_clk),
    .D(net386),
    .RESET_B(_0039_),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_1 _1455_ (.CLK(clknet_leaf_26_clk),
    .D(net370),
    .RESET_B(_0040_),
    .Q(net62));
 sky130_fd_sc_hd__dfrtp_1 _1456_ (.CLK(clknet_leaf_10_clk),
    .D(net269),
    .RESET_B(_0041_),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _1457_ (.CLK(clknet_leaf_6_clk),
    .D(net317),
    .RESET_B(_0042_),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _1458_ (.CLK(clknet_leaf_25_clk),
    .D(net305),
    .RESET_B(_0043_),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _1459_ (.CLK(clknet_leaf_25_clk),
    .D(_0262_),
    .RESET_B(_0044_),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_1 _1460_ (.CLK(clknet_leaf_12_clk),
    .D(_0263_),
    .RESET_B(_0045_),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _1461_ (.CLK(clknet_leaf_12_clk),
    .D(net303),
    .RESET_B(_0046_),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_4 _1462_ (.CLK(clknet_leaf_11_clk),
    .D(net340),
    .RESET_B(_0047_),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_1 _1463_ (.CLK(clknet_leaf_7_clk),
    .D(net395),
    .RESET_B(_0048_),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_1 _1464_ (.CLK(clknet_leaf_20_clk),
    .D(net307),
    .RESET_B(_0049_),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _1465_ (.CLK(clknet_leaf_0_clk),
    .D(net232),
    .RESET_B(_0050_),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 _1466_ (.CLK(clknet_leaf_19_clk),
    .D(net322),
    .RESET_B(_0051_),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _1467_ (.CLK(clknet_leaf_11_clk),
    .D(net142),
    .RESET_B(_0052_),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _1468_ (.CLK(clknet_leaf_25_clk),
    .D(_0271_),
    .RESET_B(_0053_),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_2 _1469_ (.CLK(clknet_leaf_8_clk),
    .D(net188),
    .RESET_B(_0054_),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _1470_ (.CLK(clknet_leaf_1_clk),
    .D(net212),
    .RESET_B(_0055_),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _1471_ (.CLK(clknet_leaf_27_clk),
    .D(net324),
    .RESET_B(_0056_),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _1472_ (.CLK(clknet_leaf_20_clk),
    .D(net146),
    .RESET_B(_0057_),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_1 _1473_ (.CLK(clknet_leaf_7_clk),
    .D(net361),
    .RESET_B(_0058_),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_1 _1474_ (.CLK(clknet_leaf_8_clk),
    .D(net348),
    .RESET_B(_0059_),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_1 _1475_ (.CLK(clknet_leaf_0_clk),
    .D(net158),
    .RESET_B(_0060_),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_1 _1476_ (.CLK(clknet_leaf_26_clk),
    .D(net174),
    .RESET_B(_0061_),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _1477_ (.CLK(clknet_leaf_26_clk),
    .D(net202),
    .RESET_B(_0062_),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_2 _1478_ (.CLK(clknet_leaf_11_clk),
    .D(net180),
    .RESET_B(_0063_),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_1 _1479_ (.CLK(clknet_leaf_11_clk),
    .D(net311),
    .RESET_B(_0064_),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _1480_ (.CLK(clknet_leaf_25_clk),
    .D(_0283_),
    .RESET_B(_0065_),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_2 _1481_ (.CLK(clknet_leaf_11_clk),
    .D(_0284_),
    .RESET_B(_0066_),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_2 _1482_ (.CLK(clknet_leaf_21_clk),
    .D(_0285_),
    .RESET_B(_0067_),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_1 _1483_ (.CLK(clknet_leaf_7_clk),
    .D(_0286_),
    .RESET_B(_0068_),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_1 _1484_ (.CLK(clknet_leaf_2_clk),
    .D(_0287_),
    .RESET_B(_0069_),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_1 _1485_ (.CLK(clknet_leaf_0_clk),
    .D(_0288_),
    .RESET_B(_0070_),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_1 _1486_ (.CLK(clknet_leaf_25_clk),
    .D(_0289_),
    .RESET_B(_0071_),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_2 _1487_ (.CLK(clknet_leaf_10_clk),
    .D(_0290_),
    .RESET_B(_0072_),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_1 _1488_ (.CLK(clknet_leaf_22_clk),
    .D(net392),
    .RESET_B(_0073_),
    .Q(\uart_tx_inst.i_data_valid ));
 sky130_fd_sc_hd__dfrtp_1 _1489_ (.CLK(clknet_leaf_23_clk),
    .D(_0292_),
    .RESET_B(_0074_),
    .Q(\uart_tx_inst.i_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1490_ (.CLK(clknet_leaf_22_clk),
    .D(net196),
    .RESET_B(_0075_),
    .Q(\uart_tx_inst.i_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1491_ (.CLK(clknet_leaf_15_clk),
    .D(_0294_),
    .RESET_B(_0076_),
    .Q(\uart_tx_inst.i_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1492_ (.CLK(clknet_leaf_19_clk),
    .D(net350),
    .RESET_B(_0077_),
    .Q(\uart_tx_inst.i_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1493_ (.CLK(clknet_leaf_21_clk),
    .D(net277),
    .RESET_B(_0078_),
    .Q(\uart_tx_inst.i_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1494_ (.CLK(clknet_leaf_20_clk),
    .D(net240),
    .RESET_B(_0079_),
    .Q(\uart_tx_inst.i_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1495_ (.CLK(clknet_leaf_21_clk),
    .D(net244),
    .RESET_B(_0080_),
    .Q(\uart_tx_inst.i_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1496_ (.CLK(clknet_leaf_19_clk),
    .D(_0299_),
    .RESET_B(_0081_),
    .Q(\uart_tx_inst.i_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1497_ (.CLK(clknet_leaf_3_clk),
    .D(_0300_),
    .RESET_B(_0082_),
    .Q(\cmd_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1498_ (.CLK(clknet_leaf_3_clk),
    .D(_0301_),
    .RESET_B(_0083_),
    .Q(\cmd_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1499_ (.CLK(clknet_leaf_3_clk),
    .D(net378),
    .RESET_B(_0084_),
    .Q(\cmd_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1500_ (.CLK(clknet_leaf_2_clk),
    .D(_0303_),
    .RESET_B(_0085_),
    .Q(\cmd_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1501_ (.CLK(clknet_leaf_24_clk),
    .D(_0304_),
    .RESET_B(_0086_),
    .Q(\cmd_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1502_ (.CLK(clknet_leaf_24_clk),
    .D(_0305_),
    .RESET_B(_0087_),
    .Q(\cmd_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1503_ (.CLK(clknet_leaf_2_clk),
    .D(_0306_),
    .RESET_B(_0088_),
    .Q(\cmd_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1504_ (.CLK(clknet_leaf_2_clk),
    .D(_0307_),
    .RESET_B(_0089_),
    .Q(\cmd_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1505_ (.CLK(clknet_leaf_27_clk),
    .D(net210),
    .RESET_B(_0090_),
    .Q(\addr_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1506_ (.CLK(clknet_leaf_5_clk),
    .D(net228),
    .RESET_B(_0091_),
    .Q(\addr_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1507_ (.CLK(clknet_leaf_11_clk),
    .D(_0310_),
    .RESET_B(_0092_),
    .Q(\addr_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1508_ (.CLK(clknet_leaf_26_clk),
    .D(net301),
    .RESET_B(_0093_),
    .Q(\addr_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1509_ (.CLK(clknet_leaf_12_clk),
    .D(net331),
    .RESET_B(_0094_),
    .Q(\addr_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1510_ (.CLK(clknet_leaf_12_clk),
    .D(net294),
    .RESET_B(_0095_),
    .Q(\addr_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1511_ (.CLK(clknet_leaf_18_clk),
    .D(_0314_),
    .RESET_B(_0096_),
    .Q(\addr_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1512_ (.CLK(clknet_leaf_20_clk),
    .D(net336),
    .RESET_B(_0097_),
    .Q(\addr_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1513_ (.CLK(clknet_leaf_17_clk),
    .D(net267),
    .RESET_B(_0098_),
    .Q(\addr_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1514_ (.CLK(clknet_leaf_0_clk),
    .D(_0317_),
    .RESET_B(_0099_),
    .Q(\addr_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1515_ (.CLK(clknet_leaf_11_clk),
    .D(net262),
    .RESET_B(_0100_),
    .Q(\addr_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1516_ (.CLK(clknet_leaf_9_clk),
    .D(_0319_),
    .RESET_B(_0101_),
    .Q(\addr_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1517_ (.CLK(clknet_leaf_26_clk),
    .D(_0320_),
    .RESET_B(_0102_),
    .Q(\addr_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1518_ (.CLK(clknet_leaf_11_clk),
    .D(_0321_),
    .RESET_B(_0103_),
    .Q(\addr_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1519_ (.CLK(clknet_leaf_1_clk),
    .D(_0322_),
    .RESET_B(_0104_),
    .Q(\addr_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1520_ (.CLK(clknet_leaf_0_clk),
    .D(net280),
    .RESET_B(_0105_),
    .Q(\addr_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1521_ (.CLK(clknet_leaf_21_clk),
    .D(_0324_),
    .RESET_B(_0106_),
    .Q(\addr_reg[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1522_ (.CLK(clknet_leaf_5_clk),
    .D(_0325_),
    .RESET_B(_0107_),
    .Q(\addr_reg[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1523_ (.CLK(clknet_leaf_15_clk),
    .D(_0326_),
    .RESET_B(_0108_),
    .Q(\addr_reg[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1524_ (.CLK(clknet_leaf_5_clk),
    .D(_0327_),
    .RESET_B(_0109_),
    .Q(\addr_reg[19] ));
 sky130_fd_sc_hd__dfrtp_1 _1525_ (.CLK(clknet_leaf_12_clk),
    .D(net265),
    .RESET_B(_0110_),
    .Q(\addr_reg[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1526_ (.CLK(clknet_leaf_19_clk),
    .D(net222),
    .RESET_B(_0111_),
    .Q(\addr_reg[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1527_ (.CLK(clknet_leaf_19_clk),
    .D(net298),
    .RESET_B(_0112_),
    .Q(\addr_reg[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1528_ (.CLK(clknet_leaf_14_clk),
    .D(_0331_),
    .RESET_B(_0113_),
    .Q(\addr_reg[23] ));
 sky130_fd_sc_hd__dfrtp_1 _1529_ (.CLK(clknet_leaf_10_clk),
    .D(_0332_),
    .RESET_B(_0114_),
    .Q(\addr_reg[24] ));
 sky130_fd_sc_hd__dfrtp_1 _1530_ (.CLK(clknet_leaf_5_clk),
    .D(net258),
    .RESET_B(_0115_),
    .Q(\addr_reg[25] ));
 sky130_fd_sc_hd__dfrtp_1 _1531_ (.CLK(clknet_leaf_10_clk),
    .D(_0334_),
    .RESET_B(_0116_),
    .Q(\addr_reg[26] ));
 sky130_fd_sc_hd__dfrtp_1 _1532_ (.CLK(clknet_leaf_10_clk),
    .D(net194),
    .RESET_B(_0117_),
    .Q(\addr_reg[27] ));
 sky130_fd_sc_hd__dfrtp_1 _1533_ (.CLK(clknet_leaf_26_clk),
    .D(net314),
    .RESET_B(_0118_),
    .Q(\addr_reg[28] ));
 sky130_fd_sc_hd__dfrtp_1 _1534_ (.CLK(clknet_leaf_11_clk),
    .D(_0337_),
    .RESET_B(_0119_),
    .Q(\addr_reg[29] ));
 sky130_fd_sc_hd__dfrtp_1 _1535_ (.CLK(clknet_leaf_0_clk),
    .D(_0338_),
    .RESET_B(_0120_),
    .Q(\addr_reg[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1536_ (.CLK(clknet_leaf_0_clk),
    .D(_0339_),
    .RESET_B(_0121_),
    .Q(\addr_reg[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1537_ (.CLK(clknet_leaf_10_clk),
    .D(net248),
    .RESET_B(_0122_),
    .Q(\data_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1538_ (.CLK(clknet_leaf_6_clk),
    .D(net285),
    .RESET_B(_0123_),
    .Q(\data_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1539_ (.CLK(clknet_leaf_25_clk),
    .D(net200),
    .RESET_B(_0124_),
    .Q(\data_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1540_ (.CLK(clknet_leaf_25_clk),
    .D(_0343_),
    .RESET_B(_0125_),
    .Q(\data_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1541_ (.CLK(clknet_leaf_12_clk),
    .D(_0344_),
    .RESET_B(_0126_),
    .Q(\data_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1542_ (.CLK(clknet_leaf_12_clk),
    .D(net290),
    .RESET_B(_0127_),
    .Q(\data_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1543_ (.CLK(clknet_leaf_11_clk),
    .D(net246),
    .RESET_B(_0128_),
    .Q(\data_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1544_ (.CLK(clknet_leaf_11_clk),
    .D(_0347_),
    .RESET_B(_0129_),
    .Q(\data_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1545_ (.CLK(clknet_leaf_20_clk),
    .D(_0348_),
    .RESET_B(_0130_),
    .Q(\data_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1546_ (.CLK(clknet_leaf_0_clk),
    .D(net226),
    .RESET_B(_0131_),
    .Q(\data_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1547_ (.CLK(clknet_leaf_19_clk),
    .D(net292),
    .RESET_B(_0132_),
    .Q(\data_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1548_ (.CLK(clknet_leaf_10_clk),
    .D(net220),
    .RESET_B(_0133_),
    .Q(\data_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1549_ (.CLK(clknet_leaf_25_clk),
    .D(_0352_),
    .RESET_B(_0134_),
    .Q(\data_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1550_ (.CLK(clknet_leaf_9_clk),
    .D(net309),
    .RESET_B(_0135_),
    .Q(\data_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1551_ (.CLK(clknet_leaf_1_clk),
    .D(net218),
    .RESET_B(_0136_),
    .Q(\data_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1552_ (.CLK(clknet_leaf_0_clk),
    .D(net283),
    .RESET_B(_0137_),
    .Q(\data_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1553_ (.CLK(clknet_leaf_21_clk),
    .D(net254),
    .RESET_B(_0138_),
    .Q(\data_reg[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1554_ (.CLK(clknet_leaf_5_clk),
    .D(_0357_),
    .RESET_B(_0139_),
    .Q(\data_reg[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1555_ (.CLK(clknet_leaf_9_clk),
    .D(_0358_),
    .RESET_B(_0140_),
    .Q(\data_reg[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1556_ (.CLK(clknet_leaf_0_clk),
    .D(net230),
    .RESET_B(_0141_),
    .Q(\data_reg[19] ));
 sky130_fd_sc_hd__dfrtp_1 _1557_ (.CLK(clknet_leaf_26_clk),
    .D(net273),
    .RESET_B(_0142_),
    .Q(\data_reg[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1558_ (.CLK(clknet_leaf_26_clk),
    .D(net251),
    .RESET_B(_0143_),
    .Q(\data_reg[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1559_ (.CLK(clknet_leaf_14_clk),
    .D(_0362_),
    .RESET_B(_0144_),
    .Q(\data_reg[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1560_ (.CLK(clknet_leaf_14_clk),
    .D(_0363_),
    .RESET_B(_0145_),
    .Q(\data_reg[23] ));
 sky130_fd_sc_hd__dfrtp_1 _1561_ (.CLK(clknet_leaf_24_clk),
    .D(_0364_),
    .RESET_B(_0146_),
    .Q(\byte_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1562_ (.CLK(clknet_leaf_24_clk),
    .D(_0365_),
    .RESET_B(_0147_),
    .Q(\byte_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1563_ (.CLK(clknet_leaf_21_clk),
    .D(_0366_),
    .RESET_B(_0148_),
    .Q(\byte_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1564_ (.CLK(clknet_leaf_25_clk),
    .D(_0367_),
    .RESET_B(_0149_),
    .Q(\byte_count[3] ));
 sky130_fd_sc_hd__dfstp_1 _1565_ (.CLK(clknet_leaf_18_clk),
    .D(net2),
    .SET_B(_0150_),
    .Q(\uart_rx_inst.rx_sync_1 ));
 sky130_fd_sc_hd__dfrtp_1 _1566_ (.CLK(clknet_leaf_9_clk),
    .D(_0001_),
    .RESET_B(_0151_),
    .Q(\uart_rx_inst.receiving ));
 sky130_fd_sc_hd__dfrtp_2 _1567_ (.CLK(clknet_leaf_7_clk),
    .D(_0368_),
    .RESET_B(_0152_),
    .Q(\uart_rx_inst.clock_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1568_ (.CLK(clknet_leaf_6_clk),
    .D(net464),
    .RESET_B(_0153_),
    .Q(\uart_rx_inst.clock_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1569_ (.CLK(clknet_leaf_6_clk),
    .D(net439),
    .RESET_B(_0154_),
    .Q(\uart_rx_inst.clock_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1570_ (.CLK(clknet_leaf_6_clk),
    .D(net443),
    .RESET_B(_0155_),
    .Q(\uart_rx_inst.clock_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1571_ (.CLK(clknet_leaf_9_clk),
    .D(_0372_),
    .RESET_B(_0156_),
    .Q(\uart_rx_inst.clock_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1572_ (.CLK(clknet_leaf_9_clk),
    .D(net403),
    .RESET_B(_0157_),
    .Q(\uart_rx_inst.clock_count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1573_ (.CLK(clknet_leaf_9_clk),
    .D(net459),
    .RESET_B(_0158_),
    .Q(\uart_rx_inst.clock_count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1574_ (.CLK(clknet_leaf_9_clk),
    .D(_0375_),
    .RESET_B(_0159_),
    .Q(\uart_rx_inst.clock_count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1575_ (.CLK(clknet_leaf_8_clk),
    .D(net417),
    .RESET_B(_0160_),
    .Q(\uart_rx_inst.clock_count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1576_ (.CLK(clknet_leaf_8_clk),
    .D(net425),
    .RESET_B(_0161_),
    .Q(\uart_rx_inst.clock_count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1577_ (.CLK(clknet_leaf_8_clk),
    .D(net470),
    .RESET_B(_0162_),
    .Q(\uart_rx_inst.clock_count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1578_ (.CLK(clknet_leaf_8_clk),
    .D(net381),
    .RESET_B(_0163_),
    .Q(\uart_rx_inst.clock_count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1579_ (.CLK(clknet_leaf_7_clk),
    .D(net437),
    .RESET_B(_0164_),
    .Q(\uart_rx_inst.clock_count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1580_ (.CLK(clknet_leaf_8_clk),
    .D(net383),
    .RESET_B(_0165_),
    .Q(\uart_rx_inst.clock_count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1581_ (.CLK(clknet_leaf_7_clk),
    .D(net451),
    .RESET_B(_0166_),
    .Q(\uart_rx_inst.clock_count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1582_ (.CLK(clknet_leaf_7_clk),
    .D(_0383_),
    .RESET_B(_0167_),
    .Q(\uart_rx_inst.clock_count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1583_ (.CLK(clknet_leaf_6_clk),
    .D(_0384_),
    .RESET_B(_0168_),
    .Q(\uart_rx_inst.bit_index[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1584_ (.CLK(clknet_leaf_4_clk),
    .D(_0385_),
    .RESET_B(_0169_),
    .Q(\uart_rx_inst.bit_index[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1585_ (.CLK(clknet_leaf_5_clk),
    .D(_0386_),
    .RESET_B(_0170_),
    .Q(\uart_rx_inst.bit_index[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1586_ (.CLK(clknet_leaf_5_clk),
    .D(_0387_),
    .RESET_B(_0171_),
    .Q(\uart_rx_inst.bit_index[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1587_ (.CLK(clknet_leaf_3_clk),
    .D(net176),
    .RESET_B(_0172_),
    .Q(\uart_rx_inst.o_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1588_ (.CLK(clknet_leaf_3_clk),
    .D(net346),
    .RESET_B(_0173_),
    .Q(\uart_rx_inst.o_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1589_ (.CLK(clknet_leaf_9_clk),
    .D(net152),
    .RESET_B(_0174_),
    .Q(\uart_rx_inst.o_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1590_ (.CLK(clknet_leaf_3_clk),
    .D(net344),
    .RESET_B(_0175_),
    .Q(\uart_rx_inst.o_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1591_ (.CLK(clknet_leaf_2_clk),
    .D(net334),
    .RESET_B(_0176_),
    .Q(\uart_rx_inst.o_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1592_ (.CLK(clknet_leaf_1_clk),
    .D(net138),
    .RESET_B(_0177_),
    .Q(\uart_rx_inst.o_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1593_ (.CLK(clknet_leaf_2_clk),
    .D(net140),
    .RESET_B(_0178_),
    .Q(\uart_rx_inst.o_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1594_ (.CLK(clknet_leaf_4_clk),
    .D(net275),
    .RESET_B(_0179_),
    .Q(\uart_rx_inst.o_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1595_ (.CLK(clknet_leaf_2_clk),
    .D(net333),
    .RESET_B(_0180_),
    .Q(\uart_rx_inst.o_data_valid ));
 sky130_fd_sc_hd__dfrtp_1 _1596_ (.CLK(clknet_leaf_15_clk),
    .D(net144),
    .RESET_B(_0181_),
    .Q(\uart_tx_inst.shift_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1597_ (.CLK(clknet_leaf_22_clk),
    .D(net184),
    .RESET_B(_0182_),
    .Q(\uart_tx_inst.shift_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1598_ (.CLK(clknet_leaf_15_clk),
    .D(net271),
    .RESET_B(_0183_),
    .Q(\uart_tx_inst.shift_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1599_ (.CLK(clknet_leaf_18_clk),
    .D(net168),
    .RESET_B(_0184_),
    .Q(\uart_tx_inst.shift_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1600_ (.CLK(clknet_leaf_21_clk),
    .D(net260),
    .RESET_B(_0185_),
    .Q(\uart_tx_inst.shift_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1601_ (.CLK(clknet_leaf_20_clk),
    .D(net198),
    .RESET_B(_0186_),
    .Q(\uart_tx_inst.shift_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1602_ (.CLK(clknet_leaf_22_clk),
    .D(net156),
    .RESET_B(_0187_),
    .Q(\uart_tx_inst.shift_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1603_ (.CLK(clknet_leaf_18_clk),
    .D(net150),
    .RESET_B(_0188_),
    .Q(\uart_tx_inst.shift_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1604_ (.CLK(clknet_leaf_18_clk),
    .D(net148),
    .RESET_B(_0189_),
    .Q(\uart_tx_inst.shift_reg[9] ));
 sky130_fd_sc_hd__dfstp_1 _1605_ (.CLK(clknet_leaf_25_clk),
    .D(net136),
    .SET_B(_0190_),
    .Q(\uart_rx_inst.rx_sync_2 ));
 sky130_fd_sc_hd__dfrtp_4 _1606_ (.CLK(clknet_leaf_16_clk),
    .D(net357),
    .RESET_B(_0191_),
    .Q(\uart_tx_inst.transmitting ));
 sky130_fd_sc_hd__dfstp_1 _1607_ (.CLK(clknet_leaf_16_clk),
    .D(net467),
    .SET_B(_0192_),
    .Q(net37));
 sky130_fd_sc_hd__dfrtp_2 _1608_ (.CLK(clknet_leaf_14_clk),
    .D(net486),
    .RESET_B(_0193_),
    .Q(\uart_tx_inst.clock_count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1609_ (.CLK(clknet_leaf_14_clk),
    .D(net457),
    .RESET_B(_0194_),
    .Q(\uart_tx_inst.clock_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1610_ (.CLK(clknet_leaf_14_clk),
    .D(net420),
    .RESET_B(_0195_),
    .Q(\uart_tx_inst.clock_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1611_ (.CLK(clknet_leaf_13_clk),
    .D(net406),
    .RESET_B(_0196_),
    .Q(\uart_tx_inst.clock_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1612_ (.CLK(clknet_leaf_12_clk),
    .D(net455),
    .RESET_B(_0197_),
    .Q(\uart_tx_inst.clock_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1613_ (.CLK(clknet_leaf_13_clk),
    .D(_0411_),
    .RESET_B(_0198_),
    .Q(\uart_tx_inst.clock_count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1614_ (.CLK(clknet_leaf_13_clk),
    .D(net445),
    .RESET_B(_0199_),
    .Q(\uart_tx_inst.clock_count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1615_ (.CLK(clknet_leaf_13_clk),
    .D(_0413_),
    .RESET_B(_0200_),
    .Q(\uart_tx_inst.clock_count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1616_ (.CLK(clknet_leaf_17_clk),
    .D(net493),
    .RESET_B(_0201_),
    .Q(\uart_tx_inst.clock_count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1617_ (.CLK(clknet_leaf_17_clk),
    .D(net474),
    .RESET_B(_0202_),
    .Q(\uart_tx_inst.clock_count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1618_ (.CLK(clknet_leaf_16_clk),
    .D(net410),
    .RESET_B(_0203_),
    .Q(\uart_tx_inst.clock_count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1619_ (.CLK(clknet_leaf_17_clk),
    .D(net363),
    .RESET_B(_0204_),
    .Q(\uart_tx_inst.clock_count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1620_ (.CLK(clknet_leaf_14_clk),
    .D(net432),
    .RESET_B(_0205_),
    .Q(\uart_tx_inst.clock_count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1621_ (.CLK(clknet_leaf_16_clk),
    .D(_0419_),
    .RESET_B(_0206_),
    .Q(\uart_tx_inst.clock_count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1622_ (.CLK(clknet_leaf_14_clk),
    .D(net489),
    .RESET_B(_0207_),
    .Q(\uart_tx_inst.clock_count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1623_ (.CLK(clknet_leaf_14_clk),
    .D(net478),
    .RESET_B(_0208_),
    .Q(\uart_tx_inst.clock_count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1624_ (.CLK(clknet_leaf_18_clk),
    .D(_0422_),
    .RESET_B(_0209_),
    .Q(\uart_tx_inst.bit_index[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1625_ (.CLK(clknet_leaf_16_clk),
    .D(net453),
    .RESET_B(_0210_),
    .Q(\uart_tx_inst.bit_index[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1626_ (.CLK(clknet_leaf_17_clk),
    .D(net428),
    .RESET_B(_0211_),
    .Q(\uart_tx_inst.bit_index[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1627_ (.CLK(clknet_leaf_17_clk),
    .D(net449),
    .RESET_B(_0212_),
    .Q(\uart_tx_inst.bit_index[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1628_ (.CLK(clknet_leaf_2_clk),
    .D(net327),
    .RESET_B(_0213_),
    .Q(\uart_rx_inst.shift_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1629_ (.CLK(clknet_leaf_3_clk),
    .D(_0427_),
    .RESET_B(_0214_),
    .Q(\uart_rx_inst.shift_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1630_ (.CLK(clknet_leaf_3_clk),
    .D(net430),
    .RESET_B(_0215_),
    .Q(\uart_rx_inst.shift_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1631_ (.CLK(clknet_leaf_3_clk),
    .D(_0429_),
    .RESET_B(_0216_),
    .Q(\uart_rx_inst.shift_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1632_ (.CLK(clknet_leaf_2_clk),
    .D(net160),
    .RESET_B(_0217_),
    .Q(\uart_rx_inst.shift_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1633_ (.CLK(clknet_leaf_4_clk),
    .D(net166),
    .RESET_B(_0218_),
    .Q(\uart_rx_inst.shift_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1634_ (.CLK(clknet_leaf_1_clk),
    .D(net192),
    .RESET_B(_0219_),
    .Q(\uart_rx_inst.shift_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1635_ (.CLK(clknet_leaf_4_clk),
    .D(_0433_),
    .RESET_B(_0220_),
    .Q(\uart_rx_inst.shift_reg[7] ));
 sky130_fd_sc_hd__clkbuf_2 _1636_ (.A(net70),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__buf_6 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__buf_6 fanout106 (.A(_0468_),
    .X(net106));
 sky130_fd_sc_hd__buf_6 fanout107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__buf_6 fanout108 (.A(_0462_),
    .X(net108));
 sky130_fd_sc_hd__buf_6 fanout109 (.A(_0437_),
    .X(net109));
 sky130_fd_sc_hd__buf_8 fanout110 (.A(_0677_),
    .X(net110));
 sky130_fd_sc_hd__buf_4 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_8 fanout112 (.A(_0675_),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__buf_4 fanout114 (.A(_0675_),
    .X(net114));
 sky130_fd_sc_hd__buf_4 fanout115 (.A(net308),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_8 fanout116 (.A(net215),
    .X(net116));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__buf_4 fanout118 (.A(net229),
    .X(net118));
 sky130_fd_sc_hd__buf_8 fanout119 (.A(net135),
    .X(net119));
 sky130_fd_sc_hd__buf_8 fanout120 (.A(net135),
    .X(net120));
 sky130_fd_sc_hd__buf_8 fanout121 (.A(net135),
    .X(net121));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net135),
    .X(net122));
 sky130_fd_sc_hd__buf_8 fanout123 (.A(net126),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_8 fanout124 (.A(net126),
    .X(net124));
 sky130_fd_sc_hd__buf_8 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_8 fanout126 (.A(net135),
    .X(net126));
 sky130_fd_sc_hd__buf_8 fanout127 (.A(net135),
    .X(net127));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net135),
    .X(net128));
 sky130_fd_sc_hd__buf_8 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__buf_6 fanout130 (.A(net135),
    .X(net130));
 sky130_fd_sc_hd__buf_6 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_6 fanout132 (.A(net134),
    .X(net132));
 sky130_fd_sc_hd__buf_8 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_8 fanout135 (.A(net3),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net499),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\data_reg[16] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\addr_reg[15] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_0242_),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net38),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_0227_),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\uart_tx_inst.i_data[5] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0297_),
    .X(net240));
 sky130_fd_sc_hd__buf_1 hold106 (.A(\uart_tx_inst.o_ready ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0649_),
    .X(net242));
 sky130_fd_sc_hd__buf_2 hold108 (.A(_0442_),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0298_),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0275_),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\data_reg[6] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0346_),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\data_reg[0] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_0340_),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 hold114 (.A(net517),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_2 hold115 (.A(_0680_),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_0361_),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_2 hold117 (.A(net514),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_0685_),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0356_),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\uart_tx_inst.shift_reg[9] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\uart_tx_inst.i_data[7] ),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_2 hold121 (.A(net508),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0700_),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0333_),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\uart_tx_inst.shift_reg[5] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_0400_),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\addr_reg[10] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_0318_),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 hold128 (.A(net515),
    .X(net263));
 sky130_fd_sc_hd__buf_1 hold129 (.A(_0681_),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0404_),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_0328_),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\addr_reg[8] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_0316_),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net71),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0259_),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net281),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_0398_),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\data_reg[20] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_0360_),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\uart_rx_inst.shift_reg[7] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net255),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_0395_),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\uart_tx_inst.i_data[4] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0296_),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_2 hold143 (.A(net509),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_0688_),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_0323_),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\uart_tx_inst.i_data[2] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\data_reg[15] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0355_),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\data_reg[1] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0403_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_0341_),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(net49),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0228_),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\uart_tx_inst.i_data[0] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\data_reg[5] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_0345_),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\data_reg[10] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_0350_),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\addr_reg[5] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_0313_),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\uart_rx_inst.shift_reg[2] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(net68),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_0235_),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 hold162 (.A(net523),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_0330_),
    .X(net298));
 sky130_fd_sc_hd__buf_2 hold164 (.A(\uart_rx_inst.o_data_valid ),
    .X(net299));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold165 (.A(_0437_),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0311_),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(net98),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_0264_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(net93),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0390_),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0261_),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(net315),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0267_),
    .X(net307));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold173 (.A(\byte_count[3] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0353_),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\data_reg[23] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_0282_),
    .X(net311));
 sky130_fd_sc_hd__buf_2 hold177 (.A(net521),
    .X(net312));
 sky130_fd_sc_hd__buf_1 hold178 (.A(_0674_),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_0336_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net318),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\data_reg[8] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(net82),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0260_),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\addr_reg[17] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(net65),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_0232_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(net72),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_0269_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(net77),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_0274_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0244_),
    .X(net154));
 sky130_fd_sc_hd__buf_2 hold190 (.A(\uart_rx_inst.bit_index[1] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_0535_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_0426_),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(net39),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_0237_),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\addr_reg[4] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_0312_),
    .X(net331));
 sky130_fd_sc_hd__buf_1 hold197 (.A(net510),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_0000_),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_0392_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\uart_rx_inst.shift_reg[5] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\uart_tx_inst.i_data[6] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\addr_reg[7] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_0315_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\addr_reg[14] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_0241_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(net99),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_0265_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(net64),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_0231_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\uart_rx_inst.shift_reg[3] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_0391_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0402_),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\uart_rx_inst.shift_reg[1] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_0389_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\data_reg[18] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_0277_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\uart_tx_inst.i_data[3] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_0295_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\addr_reg[16] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_0243_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(net67),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_0234_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\data_reg[19] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\data_reg[12] ),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_2 hold221 (.A(\uart_tx_inst.bit_index[3] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_0002_),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\cmd_reg[4] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(net74),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\data_reg[17] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_0276_),
    .X(net361));
 sky130_fd_sc_hd__buf_1 hold227 (.A(\uart_tx_inst.clock_count[11] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_0417_),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\cmd_reg[0] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_0278_),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\data_reg[3] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\data_reg[4] ),
    .X(net366));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold232 (.A(\addr_reg[18] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_0245_),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\addr_reg[31] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_0258_),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\addr_reg[30] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(net96),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\cmd_reg[7] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\addr_reg[23] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\uart_rx_inst.shift_reg[4] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0250_),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(net97),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\cmd_reg[2] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_0302_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\cmd_reg[5] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\uart_rx_inst.clock_count[11] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_0379_),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\uart_rx_inst.clock_count[13] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_0381_),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\cmd_reg[1] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0430_),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(net61),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_0257_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\cmd_reg[6] ),
    .X(net387));
 sky130_fd_sc_hd__buf_1 hold253 (.A(net518),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_0256_),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_2 hold255 (.A(net513),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\uart_tx_inst.i_data_valid ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_0291_),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\cmd_reg[3] ),
    .X(net393));
 sky130_fd_sc_hd__buf_1 hold259 (.A(net516),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\addr_reg[25] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_0266_),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_4 hold261 (.A(\uart_rx_inst.receiving ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_0609_),
    .X(net397));
 sky130_fd_sc_hd__buf_1 hold263 (.A(net520),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_0251_),
    .X(net399));
 sky130_fd_sc_hd__buf_1 hold265 (.A(net511),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_0238_),
    .X(net401));
 sky130_fd_sc_hd__buf_1 hold267 (.A(\uart_rx_inst.clock_count[5] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_0373_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(net95),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0252_),
    .X(net162));
 sky130_fd_sc_hd__buf_1 hold270 (.A(\uart_tx_inst.clock_count[3] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(_0409_),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(net104),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_0226_),
    .X(net408));
 sky130_fd_sc_hd__buf_1 hold274 (.A(\uart_tx_inst.clock_count[10] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_0416_),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_2 hold276 (.A(\state[2] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(_0661_),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_2 hold278 (.A(\uart_tx_inst.bit_index[2] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(_0600_),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\addr_reg[19] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_0224_),
    .X(net415));
 sky130_fd_sc_hd__buf_1 hold281 (.A(\uart_rx_inst.clock_count[8] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_0376_),
    .X(net417));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold283 (.A(\state[0] ),
    .X(net418));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold284 (.A(\uart_tx_inst.clock_count[2] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_0408_),
    .X(net420));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold286 (.A(\addr_reg[9] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_0236_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(net88),
    .X(net423));
 sky130_fd_sc_hd__buf_1 hold289 (.A(\uart_rx_inst.clock_count[9] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_0246_),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_0377_),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_2 hold291 (.A(\uart_tx_inst.bit_index[1] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_0536_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_0424_),
    .X(net428));
 sky130_fd_sc_hd__buf_2 hold294 (.A(\uart_rx_inst.bit_index[0] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_0428_),
    .X(net430));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold296 (.A(\uart_tx_inst.clock_count[12] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_0418_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\uart_rx_inst.clock_count[15] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_0508_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_0393_),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 hold30 (.A(\uart_rx_inst.rx_sync_2 ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_0511_),
    .X(net435));
 sky130_fd_sc_hd__buf_1 hold301 (.A(\uart_rx_inst.clock_count[12] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_0380_),
    .X(net437));
 sky130_fd_sc_hd__buf_1 hold303 (.A(\uart_rx_inst.clock_count[2] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_0370_),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(net89),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(net87),
    .X(net441));
 sky130_fd_sc_hd__buf_1 hold307 (.A(\uart_rx_inst.clock_count[3] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_0371_),
    .X(net443));
 sky130_fd_sc_hd__buf_1 hold309 (.A(\uart_tx_inst.clock_count[6] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_0431_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_0412_),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\uart_tx_inst.clock_count[13] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_0543_),
    .X(net447));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold313 (.A(_0544_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_0425_),
    .X(net449));
 sky130_fd_sc_hd__buf_1 hold315 (.A(\uart_rx_inst.clock_count[14] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_0382_),
    .X(net451));
 sky130_fd_sc_hd__buf_2 hold317 (.A(\uart_tx_inst.bit_index[0] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_0423_),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_2 hold319 (.A(\uart_tx_inst.clock_count[4] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\uart_tx_inst.shift_reg[4] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_0410_),
    .X(net455));
 sky130_fd_sc_hd__buf_1 hold321 (.A(\uart_tx_inst.clock_count[1] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_0407_),
    .X(net457));
 sky130_fd_sc_hd__buf_1 hold323 (.A(\uart_rx_inst.clock_count[6] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_0374_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(net94),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(net90),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(net91),
    .X(net462));
 sky130_fd_sc_hd__buf_1 hold328 (.A(\uart_rx_inst.clock_count[1] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_0369_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_0399_),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\state[0] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(net37),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_0405_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(net92),
    .X(net468));
 sky130_fd_sc_hd__buf_1 hold334 (.A(\uart_rx_inst.clock_count[10] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(_0378_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(net70),
    .X(net471));
 sky130_fd_sc_hd__buf_1 hold337 (.A(\uart_tx_inst.clock_count[9] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_0582_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(_0415_),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\addr_reg[12] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\uart_tx_inst.clock_count[7] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(_0587_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\uart_tx_inst.clock_count[15] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(_0421_),
    .X(net478));
 sky130_fd_sc_hd__buf_1 hold344 (.A(net525),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(_0518_),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\state[0] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\uart_rx_inst.clock_count[4] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\uart_rx_inst.clock_count[3] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(_0509_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_0239_),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\uart_tx_inst.clock_count[0] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(_0406_),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\uart_tx_inst.clock_count[14] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(_0573_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_0420_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\uart_rx_inst.clock_count[0] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\uart_tx_inst.clock_count[8] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(_0583_),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_0414_),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_2 hold359 (.A(\uart_tx_inst.transmitting ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\addr_reg[6] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\uart_tx_inst.clock_count[5] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\uart_rx_inst.clock_count[4] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\uart_tx_inst.clock_count[5] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\state[1] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\uart_rx_inst.rx_sync_1 ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\uart_tx_inst.shift_reg[8] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\uart_tx_inst.shift_reg[7] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\uart_rx_inst.o_data[7] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\uart_tx_inst.shift_reg[3] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\uart_tx_inst.shift_reg[1] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_0233_),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\uart_rx_inst.o_data[0] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\uart_rx_inst.o_data[2] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\uart_rx_inst.o_data[2] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\uart_rx_inst.o_data[1] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\uart_rx_inst.o_data[7] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\uart_rx_inst.bit_index[3] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\addr_reg[11] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\addr_reg[26] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\uart_rx_inst.o_data[2] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\uart_rx_inst.o_data[0] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net272),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\uart_rx_inst.o_data[4] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\data_reg[7] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\uart_rx_inst.o_data[5] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\addr_reg[29] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\uart_rx_inst.bit_index[2] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\addr_reg[24] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\state[1] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\uart_rx_inst.o_data[3] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\uart_rx_inst.o_data[6] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\byte_count[2] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0279_),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\uart_rx_inst.clock_count[7] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\uart_rx_inst.shift_reg[6] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\uart_rx_inst.shift_reg[0] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0388_),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\addr_reg[21] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_0248_),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\data_reg[22] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0281_),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\addr_reg[13] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0240_),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\uart_tx_inst.shift_reg[2] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0397_),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_0394_),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\addr_reg[20] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0247_),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\data_reg[13] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0272_),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 hold54 (.A(net519),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0525_),
    .X(net190));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold56 (.A(_0526_),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_0432_),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\addr_reg[27] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0335_),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\data_reg[11] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\uart_tx_inst.i_data[1] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0293_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\uart_tx_inst.shift_reg[6] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0401_),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\data_reg[2] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0342_),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\data_reg[21] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_0280_),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\addr_reg[2] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0229_),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_0270_),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\addr_reg[22] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0249_),
    .X(net206));
 sky130_fd_sc_hd__buf_1 hold72 (.A(net512),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0253_),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\addr_reg[0] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_0308_),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\data_reg[14] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_0273_),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net57),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_0254_),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net288),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 hold80 (.A(\byte_count[1] ),
    .X(net215));
 sky130_fd_sc_hd__buf_2 hold81 (.A(_0686_),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0691_),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_0354_),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 hold84 (.A(net522),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_0351_),
    .X(net220));
 sky130_fd_sc_hd__buf_2 hold86 (.A(net524),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_0329_),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\addr_reg[3] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0230_),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0396_),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\data_reg[9] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_0349_),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\addr_reg[1] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0309_),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\byte_count[0] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_0359_),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net102),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0268_),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\addr_reg[28] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0255_),
    .X(net234));
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(i_start_rx),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(wb_dat_i[14]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(wb_dat_i[15]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(wb_dat_i[16]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(wb_dat_i[17]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(wb_dat_i[18]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(wb_dat_i[19]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(wb_dat_i[1]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(wb_dat_i[20]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(wb_dat_i[21]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(wb_dat_i[22]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(i_uart_rx),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(wb_dat_i[23]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(wb_dat_i[24]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(wb_dat_i[25]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(wb_dat_i[26]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(wb_dat_i[27]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(wb_dat_i[28]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(wb_dat_i[29]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(wb_dat_i[2]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(wb_dat_i[30]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(wb_dat_i[31]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input3 (.A(rst),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(wb_dat_i[3]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(wb_dat_i[4]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(wb_dat_i[5]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(wb_dat_i[6]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(wb_dat_i[7]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(wb_dat_i[8]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(wb_dat_i[9]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input4 (.A(wb_ack_i),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(wb_dat_i[0]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(wb_dat_i[10]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(wb_dat_i[11]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(wb_dat_i[12]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(wb_dat_i[13]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output100 (.A(net100),
    .X(wb_dat_o[7]));
 sky130_fd_sc_hd__buf_12 output101 (.A(net101),
    .X(wb_dat_o[8]));
 sky130_fd_sc_hd__buf_12 output102 (.A(net102),
    .X(wb_dat_o[9]));
 sky130_fd_sc_hd__buf_12 output103 (.A(net103),
    .X(wb_stb_o));
 sky130_fd_sc_hd__buf_12 output104 (.A(net104),
    .X(wb_we_o));
 sky130_fd_sc_hd__buf_12 output37 (.A(net37),
    .X(o_uart_tx));
 sky130_fd_sc_hd__buf_12 output38 (.A(net38),
    .X(wb_adr_o[0]));
 sky130_fd_sc_hd__buf_12 output39 (.A(net39),
    .X(wb_adr_o[10]));
 sky130_fd_sc_hd__buf_12 output40 (.A(net40),
    .X(wb_adr_o[11]));
 sky130_fd_sc_hd__buf_12 output41 (.A(net41),
    .X(wb_adr_o[12]));
 sky130_fd_sc_hd__buf_12 output42 (.A(net42),
    .X(wb_adr_o[13]));
 sky130_fd_sc_hd__buf_12 output43 (.A(net43),
    .X(wb_adr_o[14]));
 sky130_fd_sc_hd__buf_12 output44 (.A(net44),
    .X(wb_adr_o[15]));
 sky130_fd_sc_hd__buf_12 output45 (.A(net45),
    .X(wb_adr_o[16]));
 sky130_fd_sc_hd__buf_12 output46 (.A(net46),
    .X(wb_adr_o[17]));
 sky130_fd_sc_hd__buf_12 output47 (.A(net47),
    .X(wb_adr_o[18]));
 sky130_fd_sc_hd__buf_12 output48 (.A(net48),
    .X(wb_adr_o[19]));
 sky130_fd_sc_hd__buf_12 output49 (.A(net49),
    .X(wb_adr_o[1]));
 sky130_fd_sc_hd__buf_12 output50 (.A(net50),
    .X(wb_adr_o[20]));
 sky130_fd_sc_hd__buf_12 output51 (.A(net51),
    .X(wb_adr_o[21]));
 sky130_fd_sc_hd__buf_12 output52 (.A(net52),
    .X(wb_adr_o[22]));
 sky130_fd_sc_hd__buf_12 output53 (.A(net53),
    .X(wb_adr_o[23]));
 sky130_fd_sc_hd__buf_12 output54 (.A(net54),
    .X(wb_adr_o[24]));
 sky130_fd_sc_hd__buf_12 output55 (.A(net55),
    .X(wb_adr_o[25]));
 sky130_fd_sc_hd__buf_12 output56 (.A(net56),
    .X(wb_adr_o[26]));
 sky130_fd_sc_hd__buf_12 output57 (.A(net57),
    .X(wb_adr_o[27]));
 sky130_fd_sc_hd__buf_12 output58 (.A(net58),
    .X(wb_adr_o[28]));
 sky130_fd_sc_hd__buf_12 output59 (.A(net59),
    .X(wb_adr_o[29]));
 sky130_fd_sc_hd__buf_12 output60 (.A(net60),
    .X(wb_adr_o[2]));
 sky130_fd_sc_hd__buf_12 output61 (.A(net61),
    .X(wb_adr_o[30]));
 sky130_fd_sc_hd__buf_12 output62 (.A(net62),
    .X(wb_adr_o[31]));
 sky130_fd_sc_hd__buf_12 output63 (.A(net63),
    .X(wb_adr_o[3]));
 sky130_fd_sc_hd__buf_12 output64 (.A(net64),
    .X(wb_adr_o[4]));
 sky130_fd_sc_hd__buf_12 output65 (.A(net65),
    .X(wb_adr_o[5]));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(wb_adr_o[6]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(wb_adr_o[7]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(wb_adr_o[8]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(wb_adr_o[9]));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(wb_cyc_o));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(wb_dat_o[0]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net72),
    .X(wb_dat_o[10]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(wb_dat_o[11]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(wb_dat_o[12]));
 sky130_fd_sc_hd__buf_12 output75 (.A(net75),
    .X(wb_dat_o[13]));
 sky130_fd_sc_hd__buf_12 output76 (.A(net76),
    .X(wb_dat_o[14]));
 sky130_fd_sc_hd__buf_12 output77 (.A(net77),
    .X(wb_dat_o[15]));
 sky130_fd_sc_hd__buf_12 output78 (.A(net78),
    .X(wb_dat_o[16]));
 sky130_fd_sc_hd__buf_12 output79 (.A(net79),
    .X(wb_dat_o[17]));
 sky130_fd_sc_hd__buf_12 output80 (.A(net80),
    .X(wb_dat_o[18]));
 sky130_fd_sc_hd__buf_12 output81 (.A(net81),
    .X(wb_dat_o[19]));
 sky130_fd_sc_hd__buf_12 output82 (.A(net82),
    .X(wb_dat_o[1]));
 sky130_fd_sc_hd__buf_12 output83 (.A(net83),
    .X(wb_dat_o[20]));
 sky130_fd_sc_hd__buf_12 output84 (.A(net84),
    .X(wb_dat_o[21]));
 sky130_fd_sc_hd__buf_12 output85 (.A(net85),
    .X(wb_dat_o[22]));
 sky130_fd_sc_hd__buf_12 output86 (.A(net86),
    .X(wb_dat_o[23]));
 sky130_fd_sc_hd__buf_12 output87 (.A(net87),
    .X(wb_dat_o[24]));
 sky130_fd_sc_hd__buf_12 output88 (.A(net88),
    .X(wb_dat_o[25]));
 sky130_fd_sc_hd__buf_12 output89 (.A(net89),
    .X(wb_dat_o[26]));
 sky130_fd_sc_hd__buf_12 output90 (.A(net90),
    .X(wb_dat_o[27]));
 sky130_fd_sc_hd__buf_12 output91 (.A(net91),
    .X(wb_dat_o[28]));
 sky130_fd_sc_hd__buf_12 output92 (.A(net92),
    .X(wb_dat_o[29]));
 sky130_fd_sc_hd__buf_12 output93 (.A(net93),
    .X(wb_dat_o[2]));
 sky130_fd_sc_hd__buf_12 output94 (.A(net94),
    .X(wb_dat_o[30]));
 sky130_fd_sc_hd__buf_12 output95 (.A(net95),
    .X(wb_dat_o[31]));
 sky130_fd_sc_hd__buf_12 output96 (.A(net96),
    .X(wb_dat_o[3]));
 sky130_fd_sc_hd__buf_12 output97 (.A(net97),
    .X(wb_dat_o[4]));
 sky130_fd_sc_hd__buf_12 output98 (.A(net98),
    .X(wb_dat_o[5]));
 sky130_fd_sc_hd__buf_12 output99 (.A(net99),
    .X(wb_dat_o[6]));
endmodule

