// This is the unpowered netlist.
module core (clk,
    o_mem_write_M,
    rst,
    i_instr_ID,
    i_read_data_M,
    o_data_addr_M,
    o_pc_IF,
    o_write_data_M);
 input clk;
 output o_mem_write_M;
 input rst;
 input [31:0] i_instr_ID;
 input [31:0] i_read_data_M;
 output [31:0] o_data_addr_M;
 output [31:0] o_pc_IF;
 output [31:0] o_write_data_M;

 wire net473;
 wire net474;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ;
 wire \U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ;
 wire \U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ;
 wire \U_CONTROL_UNIT.i_branch_EX ;
 wire \U_CONTROL_UNIT.i_jump_EX ;
 wire \U_DATAPATH.U_EX_MEM.i_mem_write_EX ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[10] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[11] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[12] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[13] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[14] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[15] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[16] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[17] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[18] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[19] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[20] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[21] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[22] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[23] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[24] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[25] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[26] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[27] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[28] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[29] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[2] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[30] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[31] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[3] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[4] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[5] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[6] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[7] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[8] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[9] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_target_EX[0] ;
 wire \U_DATAPATH.U_EX_MEM.i_pc_target_EX[1] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[0] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[1] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[2] ;
 wire \U_DATAPATH.U_EX_MEM.i_rd_EX[3] ;
 wire \U_DATAPATH.U_EX_MEM.i_reg_write_EX ;
 wire \U_DATAPATH.U_EX_MEM.i_result_src_EX[0] ;
 wire \U_DATAPATH.U_EX_MEM.i_result_src_EX[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[10] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[11] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[12] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[13] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[14] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[15] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[16] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[17] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[18] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[19] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[20] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[21] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[22] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[23] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[24] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[25] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[26] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[27] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[28] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[29] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[30] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[31] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[4] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[5] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[6] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[7] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[8] ;
 wire \U_DATAPATH.U_EX_MEM.o_alu_result_M[9] ;
 wire \U_DATAPATH.U_EX_MEM.o_mem_write_M ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[10] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[11] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[12] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[13] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[14] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[15] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[16] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[17] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[18] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[19] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[20] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[21] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[22] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[23] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[24] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[25] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[26] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[27] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[28] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[29] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[30] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[31] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[4] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[5] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[6] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[7] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[8] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_plus4_M[9] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[10] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[11] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[12] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[13] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[14] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[15] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[16] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[17] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[18] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[19] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[20] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[21] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[22] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[23] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[24] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[25] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[26] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[27] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[28] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[29] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[30] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[31] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[4] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[5] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[6] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[7] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[8] ;
 wire \U_DATAPATH.U_EX_MEM.o_pc_target_M[9] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_rd_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_reg_write_M ;
 wire \U_DATAPATH.U_EX_MEM.o_result_src_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_result_src_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[0] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[10] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[11] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[12] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[13] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[14] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[15] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[16] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[17] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[18] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[19] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[1] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[20] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[21] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[22] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[23] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[24] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[25] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[26] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[27] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[28] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[29] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[2] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[30] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[31] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[3] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[4] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[5] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[6] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[7] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[8] ;
 wire \U_DATAPATH.U_EX_MEM.o_write_data_M[9] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ;
 wire \U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_pc_plus4_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[0] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[1] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_rd_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[0] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[1] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_rs1_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[0] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[10] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[11] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[12] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[13] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[14] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[15] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[16] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[17] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[18] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[19] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[1] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[20] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[21] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[22] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[23] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[24] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[25] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[26] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[27] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[28] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[29] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[2] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[30] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[31] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[3] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[4] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[5] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[6] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[7] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[8] ;
 wire \U_DATAPATH.U_ID_EX.i_rs2_ID[9] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_alu_src_EX ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_pc_EX[9] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_rs1_EX[9] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[0] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[10] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[11] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[12] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[13] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[14] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[15] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[16] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[17] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[18] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[19] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[1] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[20] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[21] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[22] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[23] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[24] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[25] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[26] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[27] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[28] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[29] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[2] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[30] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[31] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[3] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[4] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[5] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[6] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[7] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[8] ;
 wire \U_DATAPATH.U_ID_EX.o_rs2_EX[9] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[10] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[11] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[12] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[13] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[14] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[15] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[16] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[17] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[18] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[19] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[20] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[21] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[22] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[23] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[24] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[25] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[26] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[27] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[28] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[29] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[2] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[30] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[31] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[3] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[4] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[5] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[6] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[7] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[8] ;
 wire \U_DATAPATH.U_IF_ID.i_pcplus4_IF[9] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[11] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[19] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[24] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[25] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[26] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[27] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[28] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[29] ;
 wire \U_DATAPATH.U_IF_ID.o_instr_ID[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[1] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_alu_result_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[1] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_pc_target_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[10] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[11] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[12] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[13] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[14] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[15] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[16] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[17] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[18] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[19] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[1] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[20] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[21] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[22] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[23] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[24] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[25] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[26] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[27] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[28] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[29] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[2] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[30] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[31] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[3] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[4] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[5] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[6] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[7] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[8] ;
 wire \U_DATAPATH.U_MEM_WB.o_read_data_WB[9] ;
 wire \U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ;
 wire \U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ;
 wire \U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_9_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net21;
 wire net210;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net211;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net212;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net213;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net216;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net217;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net218;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net219;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net22;
 wire net220;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net221;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net222;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net223;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net235;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net236;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net237;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net238;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net239;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net24;
 wire net240;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net241;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net242;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net243;
 wire net2430;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net2308));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_3354_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net2303));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_1811_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net1999));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net2261));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net2263));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__B (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__B (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__B (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__A_N (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__B (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A1 (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__B2 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A1 (.DIODE(_1461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__S (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__A (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A1 (.DIODE(net2190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__B2 (.DIODE(_1469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A (.DIODE(net2190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__B1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__A1 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__S (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__B1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A2 (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__B2 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__B (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__B (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A1 (.DIODE(net2035));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__B2 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A1 (.DIODE(net2035));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A2 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__A (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__A (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A1 (.DIODE(_1505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__B1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__B (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__B (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A1 (.DIODE(_1518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A1 (.DIODE(net2007));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__B2 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__C_N (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A (.DIODE(net2007));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__B (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__B1_N (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__A1 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__S (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A1 (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__B2 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A1 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__S (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A1 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__B2 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A1 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__S (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A (.DIODE(net2253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__B1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A1 (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__S (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A1 (.DIODE(net2253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__B2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__B (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__B (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A1 (.DIODE(net2077));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__B2 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__B1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__A1 (.DIODE(net2077));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__A2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__S0 (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__S1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A (.DIODE(net2167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__A1 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__S (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__B (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A1 (.DIODE(net2167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__B2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__B (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__B (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__B2 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__B (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A1 (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__S (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__A (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A1 (.DIODE(_1613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__B1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A1 (.DIODE(net2045));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A2 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A2 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A1 (.DIODE(net2045));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__B (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__B (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A1 (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__B2 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__B1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A1 (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__S (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A_N (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A1 (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__B1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A1 (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__S (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__A_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A1 (.DIODE(_1651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__B2 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__B1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__B (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A2 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__A2 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__A1 (.DIODE(_1664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A2 (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__B2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__B1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__B (.DIODE(net2162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A2 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A2 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__B (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__B (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A2 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__A2 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__B2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__B (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__A (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A_N (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__C (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__B (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A_N (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__B1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__B2 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__A1 (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__B2 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A1 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__S (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__A (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__B (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__B1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A2 (.DIODE(_1719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A2 (.DIODE(_1719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__B (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__B (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__A_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__B2 (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__B1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A1 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__S (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A1 (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__B2 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__B1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A1 (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__S (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A_N (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__B2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__A1 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__S (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__A (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__A (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__B1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__B (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__B (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A_N (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A1 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A1 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__S (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__A (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__A (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__B2 (.DIODE(\U_DATAPATH.U_MEM_WB.o_read_data_WB[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A1 (.DIODE(net2191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A2 (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__B1 (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__B2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__A (.DIODE(net2191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__B1 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__A1 (.DIODE(_1791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__S (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__A (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__A (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__A_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__B1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A0 (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A1 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__S (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A (.DIODE(net2137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A0 (.DIODE(net2332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__S (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A1 (.DIODE(net2137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__B2 (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__B (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__A1 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__S (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__B1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__A1 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__S (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__A (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A2 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A1 (.DIODE(_1831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__S (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A1 (.DIODE(net1970));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__A (.DIODE(net1970));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A0 (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A1 (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__S (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__C (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A_N (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__A_N (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__A_N (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__A2 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A_N (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__A2 (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__B2 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__A_N (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__A2 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__A_N (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A_N (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__A2 (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__B2 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__A_N (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A_N (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__A_N (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__B1 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__A_N (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A2 (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__B2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__A_N (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__A_N (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__A3 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__B2 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__A_N (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__A (.DIODE(net2162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__A (.DIODE(net2162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__S (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A1 (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__S (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__S (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__A (.DIODE(net2332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__S (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__B (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A2 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__S (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__S (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__S (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__S (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__S (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__S (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__S (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__S (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__S (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__S (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__A1_N (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__A1 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__S (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__B (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__A2 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A1 (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__A (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__A (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__S (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__B (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__S (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__S (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__S (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__S (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__S (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__S (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__S (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__S (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__A_N (.DIODE(net2210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__B (.DIODE(net2254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__A_N (.DIODE(net2258));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__B (.DIODE(net2170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__B (.DIODE(net2170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__C_N (.DIODE(net2258));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__S0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__S1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__S0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__S1 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__S1 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__S1 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__S1 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__S1 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__S1 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__S0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__S1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__S (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__S1 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__S0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__S1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__S (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__S0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__S (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__S1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__S0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__S (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__S (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__S1 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__S1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__S1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__S0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__S1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__S (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__B (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__B (.DIODE(net2191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__B (.DIODE(net2137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__B (.DIODE(net1970));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__B (.DIODE(net2007));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__B (.DIODE(net2045));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__B (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__B (.DIODE(net2190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__B (.DIODE(net2035));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__B (.DIODE(net2253));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__B (.DIODE(net2077));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__B (.DIODE(net2167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__S1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__S1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__S1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__S1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__S1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__S1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__S0 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__S (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__S1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__S1 (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__S1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__S1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__S (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__S1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__S1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__S1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__S0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__S1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__S1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__S0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__S1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__S1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__S1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__S1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__S0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__S0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__S1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__S (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__S (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__B (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A (.DIODE(net2254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A (.DIODE(net2210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A1 (.DIODE(net2258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__S (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__C_N (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__A1 (.DIODE(net2170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__S (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__C_N (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A (.DIODE(net2145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__B1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__B1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__B1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A (.DIODE(net2109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__B1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A (.DIODE(net2188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A (.DIODE(net1878));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A (.DIODE(net2175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A (.DIODE(net1971));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A (.DIODE(net2048));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A (.DIODE(net2090));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__B1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A1 (.DIODE(_1832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__B (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A1 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A (.DIODE(net2145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__C (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__A (.DIODE(net2210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__B (.DIODE(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A (.DIODE(net2170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__B (.DIODE(net2258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A_N (.DIODE(net2145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A (.DIODE(net2145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A2 (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__B (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__C_N (.DIODE(net2258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A (.DIODE(net2258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__C_N (.DIODE(net2170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A (.DIODE(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__C_N (.DIODE(net2170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__B (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A2 (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A1 (.DIODE(net2145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A (.DIODE(net2210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__B (.DIODE(net2254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A (.DIODE(net1989));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__B (.DIODE(net2170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A2 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__C (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__C (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__C (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__C (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__C (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__C (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__C (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__C (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__C (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__C (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__C (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__C (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__C (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__C (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__C (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__C (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__C (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__C (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__C (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__C (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__C (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__C (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__C (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__C (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__C (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__C (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__C (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__C (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__C (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__C (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__C (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__C (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__C (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__C (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__C (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__B (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__A1 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__A2 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__A3 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__S0 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__S1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A0 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A1 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A0 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A1 (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A2 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A3 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__S0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__S1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A0 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__S (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A0 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__S (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A0 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A1 (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__S (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A0 (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A1 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__S (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A0 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__S (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A0 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__S (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A0 (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__S (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__S (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A0 (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A1 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__S (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__S (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__S (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__S (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__B1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A_N (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__B1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__B2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__B (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__C1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A0 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A1 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__S (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__A0 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__A1 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__A2 (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__A3 (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__S1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A0 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A3 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__S0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A0 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A1 (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A2 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A3 (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__S0 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A1 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__S (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__C (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__S (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__B1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__S (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A2 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__S0 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__S1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A1 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A2 (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A3 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A0 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A1 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A0 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A2 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A3 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A0 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__S (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__S (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__S (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__S (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__A2 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__A3 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A1 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A2 (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A3 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__S (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__S (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__S (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__S (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__B (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__B1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A2 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A2 (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__B2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__B1_N (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__C1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A0 (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A1 (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A3 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__S1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A0 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A1 (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A3 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A0 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A1 (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A2 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A3 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__S1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__B (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__B1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__B1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__B2 (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A1 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A2 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A3 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__S1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A0 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A1 (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A2 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A3 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__S1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__S (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__S (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__C1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__B (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__A2 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__S1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__S (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__S1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__B1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A3 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A2 (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__C1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__A (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__B1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A2 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A3 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5913__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5913__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__C1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__A (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__S (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__B1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__B1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A2 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A1 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A2 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A3 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__C1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__B1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A1 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A2 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A3 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__S0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__S1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A1_N (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__B1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__B (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__A (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__B1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__A2 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A1 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A2 (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A3 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__S0 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__C1 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__B1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__A (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__A (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__A (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__A1 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__A2 (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__A3 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__B1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__6004__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6004__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__C1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__B1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__A2 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A0 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A1 (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A2 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A3 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__C1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__A (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__A (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A0 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A1 (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A2 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A3 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__S0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__S1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__C1 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__B1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__B1 (.DIODE(_3075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__B1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__A (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__A (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__B1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__A2 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__B1 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A0 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A2 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A3 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__C1 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__C1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A0 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A1 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A2 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__B1 (.DIODE(_2770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A1_N (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__B1 (.DIODE(_3114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__B1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A0 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A1 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__S (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__A1 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__B1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A2 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__A2 (.DIODE(_2770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__B1 (.DIODE(_3132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__B1_N (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__C1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__A (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__B1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A1 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A2 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__S0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__S1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__C1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__B2 (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__A (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__B1 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__A (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__A (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A0 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A2 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__S0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__S1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__C1 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__C1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__B2 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A2 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__B1 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__B1 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__A (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__A (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__A0 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__A3 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__S1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__C1 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__C1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__B2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__B1 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__B1_N (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__C1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__A (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__A (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A0 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A1 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A2 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A3 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__S0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__S1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__S (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__A1 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__C1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__B2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__B2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__C1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__A (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__A (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__A0 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__A2 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__A3 (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__S (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__C1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__B2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__B1 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__A1 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__C1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__B (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__A (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__A (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A3 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__B1 (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A0 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A1 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A2 (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A3 (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__C1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__B1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__A (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__A (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__B1 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__C1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__A0 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__A1 (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__A2 (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__A3 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6236__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6236__C1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__C1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__A (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__A (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A0 (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A1 (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A3 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__B1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__B1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__A0 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__A1 (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__A3 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__S0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__S1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__C1 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__C1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A2 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__B2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__B1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6280__A (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6281__A (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A0 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A3 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__S0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__S1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__C1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__A2 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__C1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__C1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__A (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__A (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A0 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A3 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__S1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__A1 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__C1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__A (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__A (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6318__A (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A0 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A1 (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A3 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__B2 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__B2 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__C1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__A (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__A (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__A (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__B1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__A0 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__A2 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__A3 (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__B2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__B2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__B1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__A (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__B1_N (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A0 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A1 (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A2 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A3 (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__A1 (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__B1 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__B1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__A (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A0 (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A2 (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A3 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__A1_N (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6378__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__B1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__A (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__A (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A0 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A1 (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A2 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A3 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__C1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__C1 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__B1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__B1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__B (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__B (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__B (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__C1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A1 (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A2 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A3 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__S0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__S1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__S (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__B1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__B1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__B2 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__C1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__B (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__B1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__B (.DIODE(net2161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__B (.DIODE(net2298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__B (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__B (.DIODE(net2241));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__B (.DIODE(net2159));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__B1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__B (.DIODE(net2289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__B (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__B (.DIODE(net2266));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__B (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__B (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__B (.DIODE(net2293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__B (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__B (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__B (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__S (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__S (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__S (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__S (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6461__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6498__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6544__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6547__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__A (.DIODE(net1989));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A1 (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__C_N (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__A1 (.DIODE(net2048));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__A2 (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__C (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__A1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__B (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__B (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__A1 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A1 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__C (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__A1 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__A3 (.DIODE(_3485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__A1 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__A1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__A1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__A1 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__C (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6845__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6846__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6846__A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__A3 (.DIODE(_3519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__A1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__A1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6862__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6862__A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__A3 (.DIODE(_3519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__A1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6881__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6881__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__A1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__A1 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__A (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__A (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__B2 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6924__A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6924__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6926__A1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__6926__A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__A1 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__A1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__B2 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6948__A1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6948__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6958__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6962__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6962__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6964__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__6964__A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__A1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6968__A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6968__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__A1 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__B (.DIODE(_3552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__A3 (.DIODE(_3553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__A_N (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__C (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6984__A0 (.DIODE(net2048));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__A_N (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6990__A0 (.DIODE(net2048));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__A1 (.DIODE(net2145));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__A1_N (.DIODE(net2048));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__A1 (.DIODE(net2048));
 sky130_fd_sc_hd__diode_2 ANTENNA__6998__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__7009__A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__7012__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__7016__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__7017__A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__7018__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__7019__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__7020__A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__7023__A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__7024__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__7029__A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__A (.DIODE(net2090));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__C (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__A (.DIODE(net2090));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__B (.DIODE(net1989));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__A (.DIODE(net2048));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__B (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7033__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__A (.DIODE(net1971));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__B (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__A (.DIODE(net2175));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__B (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__A (.DIODE(net1878));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__B (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__A (.DIODE(net2188));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__B (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7041__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__B (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__A (.DIODE(net2109));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__B (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7048__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__7048__B (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__B (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__A (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__B (.DIODE(net1989));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7054__B (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__B (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__C_N (.DIODE(net2090));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__A2 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__B (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7058__A1 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7058__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7059__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__7059__B (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7060__A1 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7060__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7061__A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__7061__B (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__A1 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__B (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__A1 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__7065__A (.DIODE(net2145));
 sky130_fd_sc_hd__diode_2 ANTENNA__7065__B (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__A1 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__B (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__A1 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__A (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__B (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__A1 (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__B (.DIODE(_3620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7072__B2 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__7074__A (.DIODE(net2048));
 sky130_fd_sc_hd__diode_2 ANTENNA__7074__C (.DIODE(net1989));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__A (.DIODE(net1971));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__C (.DIODE(net1989));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__A (.DIODE(net2175));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__C (.DIODE(net1989));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__A (.DIODE(net1878));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__C (.DIODE(net1989));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__A (.DIODE(net2188));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__C (.DIODE(net1989));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__C (.DIODE(net1989));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__B2 (.DIODE(net2109));
 sky130_fd_sc_hd__diode_2 ANTENNA__7082__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__B2 (.DIODE(net2181));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__7085__B2 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__A1 (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__B2 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__A1 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__A3 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7098__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7102__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7105__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__7109__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7118__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7119__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7120__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7121__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7254__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7256__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7258__A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__7259__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7260__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7261__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7262__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7263__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7264__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__7265__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__7266__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__7267__A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__7268__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7269__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7270__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7271__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7272__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7273__A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__7274__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7275__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7276__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7277__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7278__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7279__A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__7280__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7281__A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__7284__RESET_B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__7597__D (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7871__CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7872__D (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7873__D (.DIODE(_0849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7879__D (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7903__D (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7904__D (.DIODE(net2308));
 sky130_fd_sc_hd__diode_2 ANTENNA__7906__D (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7911__D (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7923__D (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7929__D (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7930__D (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8005__D (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8026__D (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8028__D (.DIODE(_1004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8030__D (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_100_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_101_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_102_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_103_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_104_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_105_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_106_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_107_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_108_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_109_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_110_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_111_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_112_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_113_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_114_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_115_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_116_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_95_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_96_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_97_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_98_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_99_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net2115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net2115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net2115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net2115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net2115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net2115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(_3474_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(_3474_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(_3553_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(_3552_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(_3519_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(_3485_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(_3485_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(_3484_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(_3484_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(_3472_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(_3472_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(_3427_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(_3427_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_A (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_A (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout311_A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout312_A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout313_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout315_A (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout316_A (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout317_A (.DIODE(_1832_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout319_A (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout321_A (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout326_A (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout332_A (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout335_A (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout336_A (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout340_A (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout342_A (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout344_A (.DIODE(_1469_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout345_A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout346_A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout349_A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout350_A (.DIODE(_2770_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout356_A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout357_A (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout358_A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout360_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout364_A (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout365_A (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout368_A (.DIODE(net2181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout369_A (.DIODE(net2181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout370_A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout371_A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout372_A (.DIODE(net2242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout373_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout374_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout375_A (.DIODE(net2242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout376_A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout377_A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout378_A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout379_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout380_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout381_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout382_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout383_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout384_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout385_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout387_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout388_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout389_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout391_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout392_A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout393_A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout394_A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout395_A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout397_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout398_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout400_A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout401_A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout402_A (.DIODE(net2351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout403_A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout404_A (.DIODE(net2351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout405_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout406_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout407_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout408_A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout409_A (.DIODE(net2334));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout410_A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout411_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout412_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout413_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout414_A (.DIODE(net2334));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout415_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout416_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout417_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout418_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout419_A (.DIODE(net2352));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout420_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout421_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout422_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout423_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout424_A (.DIODE(net2352));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout425_A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout426_A (.DIODE(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout427_A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout428_A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout429_A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout430_A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout431_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout432_A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout433_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout434_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout436_A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout437_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout438_A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout439_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout440_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout441_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout442_A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout443_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout444_A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout445_A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout446_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout447_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout448_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout449_A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout450_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout451_A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout452_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout453_A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout454_A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout455_A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout456_A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout457_A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout458_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout459_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout461_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout462_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout463_A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout464_A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout465_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout466_A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout467_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout468_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout469_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1429_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1439_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1441_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1442_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1452_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1453_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1454_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1464_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1465_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1467_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1469_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1470_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1474_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1476_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1481_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1484_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1488_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1491_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1492_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1493_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1498_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1503_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1512_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1522_A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1540_A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1554_A (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1556_A (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1557_A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1570_A (.DIODE(\U_DATAPATH.U_IF_ID.o_instr_ID[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1576_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1583_A (.DIODE(\U_DATAPATH.U_IF_ID.o_instr_ID[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1588_A (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1595_A (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1605_A (.DIODE(\U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1617_A (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1632_A (.DIODE(_1791_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1636_A (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1641_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1649_A (.DIODE(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1650_A (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1652_A (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1653_A (.DIODE(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1656_A (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1658_A (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1661_A (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1663_A (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1676_A (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1680_A (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1684_A (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1686_A (.DIODE(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1688_A (.DIODE(_1461_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1693_A (.DIODE(_1719_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1695_A (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1698_A (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1703_A (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1729_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1744_A (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1746_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1747_A (.DIODE(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1759_A (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1761_A (.DIODE(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1765_A (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1772_A (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1780_A (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1786_A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap355_A (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_output152_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_84 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _3646_ (.A(net463),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _3647_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .Y(_1400_));
 sky130_fd_sc_hd__inv_2 _3648_ (.A(net375),
    .Y(_1401_));
 sky130_fd_sc_hd__clkinv_4 _3649_ (.A(net389),
    .Y(_1402_));
 sky130_fd_sc_hd__inv_2 _3650_ (.A(net1980),
    .Y(_1403_));
 sky130_fd_sc_hd__inv_2 _3651_ (.A(net1957),
    .Y(_1404_));
 sky130_fd_sc_hd__inv_2 _3652_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .Y(_1405_));
 sky130_fd_sc_hd__inv_2 _3653_ (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ),
    .Y(_1406_));
 sky130_fd_sc_hd__inv_2 _3654_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .Y(_1407_));
 sky130_fd_sc_hd__inv_2 _3655_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .Y(_1408_));
 sky130_fd_sc_hd__inv_2 _3656_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .Y(_1409_));
 sky130_fd_sc_hd__inv_2 _3657_ (.A(net366),
    .Y(_1410_));
 sky130_fd_sc_hd__inv_2 _3658_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .Y(_1411_));
 sky130_fd_sc_hd__inv_2 _3659_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ),
    .Y(_1412_));
 sky130_fd_sc_hd__inv_2 _3660_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ),
    .Y(_1413_));
 sky130_fd_sc_hd__inv_2 _3661_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ),
    .Y(_1414_));
 sky130_fd_sc_hd__inv_2 _3662__1 (.A(clknet_leaf_50_clk),
    .Y(net477));
 sky130_fd_sc_hd__or4_1 _3663_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ),
    .C(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ),
    .D(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ),
    .X(_1415_));
 sky130_fd_sc_hd__o2bb2a_1 _3664_ (.A1_N(_1414_),
    .A2_N(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .B1(_1406_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .X(_1416_));
 sky130_fd_sc_hd__o22a_1 _3665_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .A2(_1413_),
    .B1(_1414_),
    .B2(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .X(_1417_));
 sky130_fd_sc_hd__a22oi_1 _3666_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .A2(_1412_),
    .B1(_1413_),
    .B2(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .Y(_1418_));
 sky130_fd_sc_hd__o211a_1 _3667_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .A2(_1412_),
    .B1(_1415_),
    .C1(\U_DATAPATH.U_EX_MEM.o_reg_write_M ),
    .X(_1419_));
 sky130_fd_sc_hd__o2111a_1 _3668_ (.A1(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ),
    .A2(_1411_),
    .B1(_1417_),
    .C1(_1418_),
    .D1(_1419_),
    .X(_1420_));
 sky130_fd_sc_hd__nand2_4 _3669_ (.A(_1416_),
    .B(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__nand2b_1 _3670_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .Y(_1422_));
 sky130_fd_sc_hd__o221a_1 _3671_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .A2(_1412_),
    .B1(_1414_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .C1(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__xnor2_1 _3672_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ),
    .Y(_1424_));
 sky130_fd_sc_hd__o221a_1 _3673_ (.A1(_1407_),
    .A2(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ),
    .B1(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ),
    .B2(_1409_),
    .C1(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__o211a_1 _3674_ (.A1(_1408_),
    .A2(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ),
    .B1(_1415_),
    .C1(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .X(_1426_));
 sky130_fd_sc_hd__and3_1 _3675_ (.A(_1423_),
    .B(_1425_),
    .C(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__nand2_2 _3676_ (.A(net274),
    .B(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__nor2_1 _3677_ (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(net426),
    .Y(_1429_));
 sky130_fd_sc_hd__or2_2 _3678_ (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(net426),
    .X(_1430_));
 sky130_fd_sc_hd__and2_1 _3679_ (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(net426),
    .X(_1431_));
 sky130_fd_sc_hd__and2b_1 _3680_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[25] ),
    .X(_1432_));
 sky130_fd_sc_hd__and2b_1 _3681_ (.A_N(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(net426),
    .X(_1433_));
 sky130_fd_sc_hd__a221o_2 _3682_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[25] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[25] ),
    .C1(_1432_),
    .X(_1434_));
 sky130_fd_sc_hd__mux2_1 _3683_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[25] ),
    .A1(_1434_),
    .S(net362),
    .X(_1435_));
 sky130_fd_sc_hd__a21o_2 _3684_ (.A1(_1416_),
    .A2(_1420_),
    .B1(_1427_),
    .X(_1436_));
 sky130_fd_sc_hd__or2_1 _3685_ (.A(net2365),
    .B(net271),
    .X(_1437_));
 sky130_fd_sc_hd__o221a_4 _3686_ (.A1(net2105),
    .A2(net273),
    .B1(net243),
    .B2(net348),
    .C1(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__nand2b_1 _3687_ (.A_N(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .Y(_1439_));
 sky130_fd_sc_hd__and2b_1 _3688_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .B(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .X(_1440_));
 sky130_fd_sc_hd__nand2b_1 _3689_ (.A_N(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .Y(_1441_));
 sky130_fd_sc_hd__nor4_1 _3690_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ),
    .C(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .D(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .Y(_1442_));
 sky130_fd_sc_hd__a221o_1 _3691_ (.A1(_1405_),
    .A2(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .B1(_1406_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .C1(_1440_),
    .X(_1443_));
 sky130_fd_sc_hd__nand2_1 _3692_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .Y(_1444_));
 sky130_fd_sc_hd__or2_1 _3693_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .X(_1445_));
 sky130_fd_sc_hd__a21o_1 _3694_ (.A1(_1444_),
    .A2(_1445_),
    .B1(_1442_),
    .X(_1446_));
 sky130_fd_sc_hd__o2111ai_1 _3695_ (.A1(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .A2(_1406_),
    .B1(_1439_),
    .C1(_1441_),
    .D1(\U_DATAPATH.U_EX_MEM.o_reg_write_M ),
    .Y(_1447_));
 sky130_fd_sc_hd__nor3_1 _3696_ (.A(_1443_),
    .B(_1446_),
    .C(_1447_),
    .Y(_1448_));
 sky130_fd_sc_hd__and2b_1 _3697_ (.A_N(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .X(_1449_));
 sky130_fd_sc_hd__a2bb2o_1 _3698_ (.A1_N(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .A2_N(_1408_),
    .B1(_1409_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ),
    .X(_1450_));
 sky130_fd_sc_hd__a221o_1 _3699_ (.A1(_1405_),
    .A2(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B1(_1408_),
    .B2(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ),
    .C1(_1449_),
    .X(_1451_));
 sky130_fd_sc_hd__nand2_1 _3700_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .Y(_1452_));
 sky130_fd_sc_hd__or2_1 _3701_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .X(_1453_));
 sky130_fd_sc_hd__a21o_1 _3702_ (.A1(_1452_),
    .A2(_1453_),
    .B1(_1442_),
    .X(_1454_));
 sky130_fd_sc_hd__o21ai_1 _3703_ (.A1(_1405_),
    .A2(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B1(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .Y(_1455_));
 sky130_fd_sc_hd__nor4_1 _3704_ (.A(_1450_),
    .B(_1451_),
    .C(_1454_),
    .D(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__or4_1 _3705_ (.A(_1450_),
    .B(_1451_),
    .C(_1454_),
    .D(_1455_),
    .X(_1457_));
 sky130_fd_sc_hd__nor2_1 _3706_ (.A(net346),
    .B(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hd__and2_1 _3707_ (.A(net2105),
    .B(net345),
    .X(_1459_));
 sky130_fd_sc_hd__nor2_1 _3708_ (.A(net346),
    .B(_1456_),
    .Y(_1460_));
 sky130_fd_sc_hd__a221o_2 _3709_ (.A1(_1435_),
    .A2(net269),
    .B1(net267),
    .B2(net2292),
    .C1(_1459_),
    .X(_1461_));
 sky130_fd_sc_hd__mux2_2 _3710_ (.A0(net2328),
    .A1(_1461_),
    .S(net364),
    .X(_1462_));
 sky130_fd_sc_hd__inv_2 _3711_ (.A(_1462_),
    .Y(_1463_));
 sky130_fd_sc_hd__or2_1 _3712_ (.A(_1438_),
    .B(_1462_),
    .X(_1464_));
 sky130_fd_sc_hd__nand2_1 _3713_ (.A(_1438_),
    .B(_1462_),
    .Y(_1465_));
 sky130_fd_sc_hd__and2_1 _3714_ (.A(_1464_),
    .B(_1465_),
    .X(_1466_));
 sky130_fd_sc_hd__and2b_1 _3715_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[26] ),
    .X(_1467_));
 sky130_fd_sc_hd__a221o_1 _3716_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[26] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[26] ),
    .C1(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_2 _3717_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[26] ),
    .A1(_1468_),
    .S(net362),
    .X(_1469_));
 sky130_fd_sc_hd__or2_1 _3718_ (.A(net2363),
    .B(net271),
    .X(_1470_));
 sky130_fd_sc_hd__o221a_4 _3719_ (.A1(net2190),
    .A2(net273),
    .B1(net243),
    .B2(_1469_),
    .C1(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__and2_1 _3720_ (.A(net2190),
    .B(net345),
    .X(_1472_));
 sky130_fd_sc_hd__a221o_2 _3721_ (.A1(net2313),
    .A2(net267),
    .B1(net344),
    .B2(net269),
    .C1(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__mux2_2 _3722_ (.A0(net2318),
    .A1(_1473_),
    .S(net364),
    .X(_1474_));
 sky130_fd_sc_hd__nand2_1 _3723_ (.A(net2364),
    .B(_1474_),
    .Y(_1475_));
 sky130_fd_sc_hd__or2_1 _3724_ (.A(_1471_),
    .B(_1474_),
    .X(_1476_));
 sky130_fd_sc_hd__and2_1 _3725_ (.A(_1475_),
    .B(_1476_),
    .X(_1477_));
 sky130_fd_sc_hd__and2b_1 _3726_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[24] ),
    .X(_1478_));
 sky130_fd_sc_hd__a221o_1 _3727_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[24] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[24] ),
    .C1(_1478_),
    .X(_1479_));
 sky130_fd_sc_hd__mux2_1 _3728_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[24] ),
    .A1(_1479_),
    .S(net362),
    .X(_1480_));
 sky130_fd_sc_hd__a22o_1 _3729_ (.A1(net2138),
    .A2(net267),
    .B1(net343),
    .B2(net269),
    .X(_1481_));
 sky130_fd_sc_hd__a21oi_4 _3730_ (.A1(net2016),
    .A2(net345),
    .B1(net2139),
    .Y(_1482_));
 sky130_fd_sc_hd__nand2_1 _3731_ (.A(net366),
    .B(net2151),
    .Y(_1483_));
 sky130_fd_sc_hd__o21ai_4 _3732_ (.A1(net366),
    .A2(_1482_),
    .B1(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hd__inv_2 _3733_ (.A(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__or2_1 _3734_ (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ),
    .B(net271),
    .X(_1486_));
 sky130_fd_sc_hd__o221a_4 _3735_ (.A1(net2016),
    .A2(net273),
    .B1(net243),
    .B2(net343),
    .C1(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__nand2_1 _3736_ (.A(_1484_),
    .B(_1487_),
    .Y(_1488_));
 sky130_fd_sc_hd__or2_1 _3737_ (.A(_1484_),
    .B(_1487_),
    .X(_1489_));
 sky130_fd_sc_hd__and2b_1 _3738_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[27] ),
    .X(_1490_));
 sky130_fd_sc_hd__a221o_1 _3739_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[27] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[27] ),
    .C1(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__mux2_2 _3740_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[27] ),
    .A1(_1491_),
    .S(net362),
    .X(_1492_));
 sky130_fd_sc_hd__or2_1 _3741_ (.A(net2335),
    .B(net271),
    .X(_1493_));
 sky130_fd_sc_hd__o221a_4 _3742_ (.A1(net2035),
    .A2(net273),
    .B1(net243),
    .B2(_1492_),
    .C1(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__a22o_1 _3743_ (.A1(net2282),
    .A2(net267),
    .B1(net342),
    .B2(net269),
    .X(_1495_));
 sky130_fd_sc_hd__a21oi_4 _3744_ (.A1(net2035),
    .A2(net345),
    .B1(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__nand2_1 _3745_ (.A(net366),
    .B(net2259),
    .Y(_1497_));
 sky130_fd_sc_hd__o21ai_2 _3746_ (.A1(net366),
    .A2(_1496_),
    .B1(_1497_),
    .Y(_1498_));
 sky130_fd_sc_hd__or2_1 _3747_ (.A(_1494_),
    .B(_1498_),
    .X(_1499_));
 sky130_fd_sc_hd__nand2_1 _3748_ (.A(_1494_),
    .B(_1498_),
    .Y(_1500_));
 sky130_fd_sc_hd__and2_1 _3749_ (.A(_1499_),
    .B(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__or3_1 _3750_ (.A(_1466_),
    .B(_1477_),
    .C(_1501_),
    .X(_1502_));
 sky130_fd_sc_hd__a21o_1 _3751_ (.A1(_1488_),
    .A2(_1489_),
    .B1(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__and2b_1 _3752_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[16] ),
    .X(_1504_));
 sky130_fd_sc_hd__a221o_2 _3753_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[16] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[16] ),
    .C1(_1504_),
    .X(_1505_));
 sky130_fd_sc_hd__mux2_1 _3754_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[16] ),
    .A1(_1505_),
    .S(net362),
    .X(_1506_));
 sky130_fd_sc_hd__and2_1 _3755_ (.A(net2104),
    .B(net345),
    .X(_1507_));
 sky130_fd_sc_hd__a221o_2 _3756_ (.A1(net2199),
    .A2(net267),
    .B1(net341),
    .B2(net269),
    .C1(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__nand2_1 _3757_ (.A(net364),
    .B(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__nand2_1 _3758_ (.A(net366),
    .B(net2212),
    .Y(_1510_));
 sky130_fd_sc_hd__nand2_2 _3759_ (.A(_1509_),
    .B(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__or2_1 _3760_ (.A(net2348),
    .B(net271),
    .X(_1512_));
 sky130_fd_sc_hd__o221a_4 _3761_ (.A1(net2104),
    .A2(net273),
    .B1(net243),
    .B2(_1506_),
    .C1(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__or2_1 _3762_ (.A(_1511_),
    .B(_1513_),
    .X(_1514_));
 sky130_fd_sc_hd__nand2_1 _3763_ (.A(_1511_),
    .B(net2349),
    .Y(_1515_));
 sky130_fd_sc_hd__and2_1 _3764_ (.A(_1514_),
    .B(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__and2b_1 _3765_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[17] ),
    .X(_1517_));
 sky130_fd_sc_hd__a221o_2 _3766_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[17] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[17] ),
    .C1(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__mux2_2 _3767_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[17] ),
    .A1(_1518_),
    .S(net363),
    .X(_1519_));
 sky130_fd_sc_hd__or2_1 _3768_ (.A(net2383),
    .B(net272),
    .X(_1520_));
 sky130_fd_sc_hd__o221a_4 _3769_ (.A1(net2007),
    .A2(net274),
    .B1(net244),
    .B2(_1519_),
    .C1(_1520_),
    .X(_1521_));
 sky130_fd_sc_hd__or3b_1 _3770_ (.A(net346),
    .B(_1457_),
    .C_N(net340),
    .X(_1522_));
 sky130_fd_sc_hd__nand2_1 _3771_ (.A(net2007),
    .B(net347),
    .Y(_1523_));
 sky130_fd_sc_hd__or3b_1 _3772_ (.A(net346),
    .B(_1456_),
    .C_N(net2125),
    .X(_1524_));
 sky130_fd_sc_hd__a31o_1 _3773_ (.A1(_1522_),
    .A2(_1523_),
    .A3(_1524_),
    .B1(net367),
    .X(_1525_));
 sky130_fd_sc_hd__a21bo_2 _3774_ (.A1(net366),
    .A2(net2322),
    .B1_N(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__or2_1 _3775_ (.A(_1521_),
    .B(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__xor2_1 _3776_ (.A(_1521_),
    .B(_1526_),
    .X(_1528_));
 sky130_fd_sc_hd__and2b_1 _3777_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[18] ),
    .X(_1529_));
 sky130_fd_sc_hd__a221o_1 _3778_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[18] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[18] ),
    .C1(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__mux2_1 _3779_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[18] ),
    .A1(_1530_),
    .S(net362),
    .X(_1531_));
 sky130_fd_sc_hd__or2_1 _3780_ (.A(net2360),
    .B(net271),
    .X(_1532_));
 sky130_fd_sc_hd__o221a_4 _3781_ (.A1(net1897),
    .A2(net273),
    .B1(net243),
    .B2(net339),
    .C1(_1532_),
    .X(_1533_));
 sky130_fd_sc_hd__and2_1 _3782_ (.A(net1897),
    .B(net345),
    .X(_1534_));
 sky130_fd_sc_hd__a221o_1 _3783_ (.A1(net2288),
    .A2(net267),
    .B1(_1531_),
    .B2(net269),
    .C1(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__mux2_2 _3784_ (.A0(net2235),
    .A1(_1535_),
    .S(net364),
    .X(_1536_));
 sky130_fd_sc_hd__nand2_1 _3785_ (.A(_1533_),
    .B(_1536_),
    .Y(_1537_));
 sky130_fd_sc_hd__or2_1 _3786_ (.A(_1533_),
    .B(_1536_),
    .X(_1538_));
 sky130_fd_sc_hd__nand2_1 _3787_ (.A(_1537_),
    .B(_1538_),
    .Y(_1539_));
 sky130_fd_sc_hd__inv_2 _3788_ (.A(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__and2b_1 _3789_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[19] ),
    .X(_1541_));
 sky130_fd_sc_hd__a221o_2 _3790_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[19] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[19] ),
    .C1(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__mux2_1 _3791_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[19] ),
    .A1(_1542_),
    .S(net362),
    .X(_1543_));
 sky130_fd_sc_hd__or2_1 _3792_ (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[19] ),
    .B(net271),
    .X(_1544_));
 sky130_fd_sc_hd__o221a_4 _3793_ (.A1(net2113),
    .A2(net273),
    .B1(net243),
    .B2(net338),
    .C1(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__and2_1 _3794_ (.A(net2113),
    .B(net345),
    .X(_1546_));
 sky130_fd_sc_hd__a221o_2 _3795_ (.A1(net2284),
    .A2(net267),
    .B1(net338),
    .B2(net269),
    .C1(_1546_),
    .X(_1547_));
 sky130_fd_sc_hd__mux2_2 _3796_ (.A0(net2366),
    .A1(_1547_),
    .S(net364),
    .X(_1548_));
 sky130_fd_sc_hd__or2_1 _3797_ (.A(_1545_),
    .B(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__nand2_1 _3798_ (.A(_1545_),
    .B(_1548_),
    .Y(_1550_));
 sky130_fd_sc_hd__and2_1 _3799_ (.A(_1549_),
    .B(_1550_),
    .X(_1551_));
 sky130_fd_sc_hd__or4_1 _3800_ (.A(_1516_),
    .B(_1528_),
    .C(_1540_),
    .D(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__and2b_1 _3801_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ),
    .X(_1553_));
 sky130_fd_sc_hd__a221o_2 _3802_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[30] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[30] ),
    .C1(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__mux2_1 _3803_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[30] ),
    .A1(_1554_),
    .S(net362),
    .X(_1555_));
 sky130_fd_sc_hd__or2_1 _3804_ (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ),
    .B(net271),
    .X(_1556_));
 sky130_fd_sc_hd__o221a_4 _3805_ (.A1(net2076),
    .A2(net273),
    .B1(net243),
    .B2(net337),
    .C1(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__and2_1 _3806_ (.A(net2076),
    .B(net345),
    .X(_1558_));
 sky130_fd_sc_hd__a221o_2 _3807_ (.A1(net2280),
    .A2(net267),
    .B1(_1555_),
    .B2(net269),
    .C1(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__mux2_2 _3808_ (.A0(net2386),
    .A1(_1559_),
    .S(net364),
    .X(_1560_));
 sky130_fd_sc_hd__or2_1 _3809_ (.A(_1557_),
    .B(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__nand2_1 _3810_ (.A(_1557_),
    .B(_1560_),
    .Y(_1562_));
 sky130_fd_sc_hd__and2_1 _3811_ (.A(_1561_),
    .B(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__and2b_1 _3812_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[28] ),
    .X(_1564_));
 sky130_fd_sc_hd__a221o_1 _3813_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[28] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[28] ),
    .C1(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__mux2_2 _3814_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[28] ),
    .A1(_1565_),
    .S(net362),
    .X(_1566_));
 sky130_fd_sc_hd__and2_1 _3815_ (.A(net2253),
    .B(net345),
    .X(_1567_));
 sky130_fd_sc_hd__a221o_2 _3816_ (.A1(net2262),
    .A2(net267),
    .B1(net336),
    .B2(net269),
    .C1(_1567_),
    .X(_1568_));
 sky130_fd_sc_hd__mux2_2 _3817_ (.A0(net2201),
    .A1(_1568_),
    .S(net364),
    .X(_1569_));
 sky130_fd_sc_hd__inv_2 _3818_ (.A(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__or2_1 _3819_ (.A(net2362),
    .B(net271),
    .X(_1571_));
 sky130_fd_sc_hd__o221a_4 _3820_ (.A1(net2253),
    .A2(net273),
    .B1(net243),
    .B2(net336),
    .C1(_1571_),
    .X(_1572_));
 sky130_fd_sc_hd__or2_1 _3821_ (.A(_1569_),
    .B(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__nand2_1 _3822_ (.A(_1569_),
    .B(_1572_),
    .Y(_1574_));
 sky130_fd_sc_hd__and2_1 _3823_ (.A(_1573_),
    .B(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__and2b_1 _3824_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[29] ),
    .X(_1576_));
 sky130_fd_sc_hd__a221o_1 _3825_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[29] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[29] ),
    .C1(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__mux2_2 _3826_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[29] ),
    .A1(_1577_),
    .S(net362),
    .X(_1578_));
 sky130_fd_sc_hd__or2_1 _3827_ (.A(net2347),
    .B(net271),
    .X(_1579_));
 sky130_fd_sc_hd__o221a_4 _3828_ (.A1(net2077),
    .A2(net273),
    .B1(net243),
    .B2(net335),
    .C1(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__a22o_1 _3829_ (.A1(net2148),
    .A2(net267),
    .B1(_1578_),
    .B2(net269),
    .X(_1581_));
 sky130_fd_sc_hd__a21oi_4 _3830_ (.A1(net2077),
    .A2(net345),
    .B1(_1581_),
    .Y(_1582_));
 sky130_fd_sc_hd__nand2_1 _3831_ (.A(net366),
    .B(net2323),
    .Y(_1583_));
 sky130_fd_sc_hd__o21ai_4 _3832_ (.A1(net366),
    .A2(_1582_),
    .B1(_1583_),
    .Y(_1584_));
 sky130_fd_sc_hd__inv_2 _3833_ (.A(_1584_),
    .Y(_1585_));
 sky130_fd_sc_hd__or2_1 _3834_ (.A(_1580_),
    .B(_1584_),
    .X(_1586_));
 sky130_fd_sc_hd__nand2_1 _3835_ (.A(_1580_),
    .B(_1584_),
    .Y(_1587_));
 sky130_fd_sc_hd__and2_1 _3836_ (.A(_1586_),
    .B(_1587_),
    .X(_1588_));
 sky130_fd_sc_hd__mux4_2 _3837_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[31] ),
    .A1(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[31] ),
    .A2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[31] ),
    .A3(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[31] ),
    .S0(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .S1(net426),
    .X(_1589_));
 sky130_fd_sc_hd__and2_1 _3838_ (.A(net2167),
    .B(net345),
    .X(_1590_));
 sky130_fd_sc_hd__a221o_2 _3839_ (.A1(net2269),
    .A2(net267),
    .B1(net357),
    .B2(net269),
    .C1(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__mux2_1 _3840_ (.A0(net2353),
    .A1(_1591_),
    .S(net364),
    .X(_1592_));
 sky130_fd_sc_hd__or2_1 _3841_ (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ),
    .B(_1436_),
    .X(_1593_));
 sky130_fd_sc_hd__o221a_4 _3842_ (.A1(net2167),
    .A2(net273),
    .B1(net243),
    .B2(net357),
    .C1(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__inv_2 _3843_ (.A(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hd__nand2_1 _3844_ (.A(_1592_),
    .B(_1594_),
    .Y(_1596_));
 sky130_fd_sc_hd__or2_1 _3845_ (.A(_1592_),
    .B(_1594_),
    .X(_1597_));
 sky130_fd_sc_hd__nand2_1 _3846_ (.A(_1596_),
    .B(_1597_),
    .Y(_1598_));
 sky130_fd_sc_hd__inv_2 _3847_ (.A(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__or4_1 _3848_ (.A(_1563_),
    .B(_1575_),
    .C(_1588_),
    .D(_1599_),
    .X(_1600_));
 sky130_fd_sc_hd__and2b_1 _3849_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[22] ),
    .X(_1601_));
 sky130_fd_sc_hd__a221o_1 _3850_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[22] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[22] ),
    .C1(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__mux2_1 _3851_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[22] ),
    .A1(_1602_),
    .S(net362),
    .X(_1603_));
 sky130_fd_sc_hd__or2_1 _3852_ (.A(net2393),
    .B(net271),
    .X(_1604_));
 sky130_fd_sc_hd__o221a_4 _3853_ (.A1(net2037),
    .A2(net273),
    .B1(net243),
    .B2(net334),
    .C1(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__and2_1 _3854_ (.A(net2037),
    .B(net347),
    .X(_1606_));
 sky130_fd_sc_hd__a221o_2 _3855_ (.A1(net2265),
    .A2(net268),
    .B1(_1603_),
    .B2(net270),
    .C1(_1606_),
    .X(_1607_));
 sky130_fd_sc_hd__mux2_2 _3856_ (.A0(net2304),
    .A1(_1607_),
    .S(net364),
    .X(_1608_));
 sky130_fd_sc_hd__or2_1 _3857_ (.A(_1605_),
    .B(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__nand2_1 _3858_ (.A(_1605_),
    .B(_1608_),
    .Y(_1610_));
 sky130_fd_sc_hd__and2_1 _3859_ (.A(_1609_),
    .B(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__and2b_1 _3860_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[20] ),
    .X(_1612_));
 sky130_fd_sc_hd__a221o_2 _3861_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[20] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[20] ),
    .C1(_1612_),
    .X(_1613_));
 sky130_fd_sc_hd__mux2_1 _3862_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[20] ),
    .A1(_1613_),
    .S(net362),
    .X(_1614_));
 sky130_fd_sc_hd__a22o_1 _3863_ (.A1(net2305),
    .A2(net267),
    .B1(net333),
    .B2(net269),
    .X(_1615_));
 sky130_fd_sc_hd__a21oi_4 _3864_ (.A1(net2045),
    .A2(net345),
    .B1(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hd__nand2_1 _3865_ (.A(net366),
    .B(net2325),
    .Y(_1617_));
 sky130_fd_sc_hd__o21a_1 _3866_ (.A1(net366),
    .A2(_1616_),
    .B1(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__o21ai_1 _3867_ (.A1(net366),
    .A2(_1616_),
    .B1(_1617_),
    .Y(_1619_));
 sky130_fd_sc_hd__or2_1 _3868_ (.A(net2361),
    .B(net271),
    .X(_1620_));
 sky130_fd_sc_hd__o221a_4 _3869_ (.A1(net2045),
    .A2(net273),
    .B1(net243),
    .B2(_1614_),
    .C1(_1620_),
    .X(_1621_));
 sky130_fd_sc_hd__or2_1 _3870_ (.A(_1619_),
    .B(_1621_),
    .X(_1622_));
 sky130_fd_sc_hd__nand2_1 _3871_ (.A(_1619_),
    .B(_1621_),
    .Y(_1623_));
 sky130_fd_sc_hd__and2_1 _3872_ (.A(_1622_),
    .B(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__and2b_1 _3873_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[23] ),
    .X(_1625_));
 sky130_fd_sc_hd__a221o_1 _3874_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[23] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[23] ),
    .C1(_1625_),
    .X(_1626_));
 sky130_fd_sc_hd__mux2_2 _3875_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[23] ),
    .A1(_1626_),
    .S(net362),
    .X(_1627_));
 sky130_fd_sc_hd__or2_1 _3876_ (.A(net2390),
    .B(net271),
    .X(_1628_));
 sky130_fd_sc_hd__o221a_4 _3877_ (.A1(net2092),
    .A2(net273),
    .B1(net243),
    .B2(_1627_),
    .C1(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__and2_1 _3878_ (.A(net2092),
    .B(net345),
    .X(_1630_));
 sky130_fd_sc_hd__a221o_1 _3879_ (.A1(net2283),
    .A2(net267),
    .B1(net332),
    .B2(net269),
    .C1(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__mux2_2 _3880_ (.A0(net2329),
    .A1(_1631_),
    .S(net364),
    .X(_1632_));
 sky130_fd_sc_hd__or2_1 _3881_ (.A(_1629_),
    .B(_1632_),
    .X(_1633_));
 sky130_fd_sc_hd__nand2_1 _3882_ (.A(net2391),
    .B(_1632_),
    .Y(_1634_));
 sky130_fd_sc_hd__and2_1 _3883_ (.A(_1633_),
    .B(_1634_),
    .X(_1635_));
 sky130_fd_sc_hd__and2b_1 _3884_ (.A_N(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[21] ),
    .X(_1636_));
 sky130_fd_sc_hd__a221o_2 _3885_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[21] ),
    .A2(net361),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[21] ),
    .C1(_1636_),
    .X(_1637_));
 sky130_fd_sc_hd__mux2_1 _3886_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[21] ),
    .A1(_1637_),
    .S(net363),
    .X(_1638_));
 sky130_fd_sc_hd__or2_1 _3887_ (.A(net2376),
    .B(net272),
    .X(_1639_));
 sky130_fd_sc_hd__o221a_4 _3888_ (.A1(net2099),
    .A2(net274),
    .B1(net244),
    .B2(_1638_),
    .C1(_1639_),
    .X(_1640_));
 sky130_fd_sc_hd__and2_1 _3889_ (.A(net2099),
    .B(net346),
    .X(_1641_));
 sky130_fd_sc_hd__a221o_2 _3890_ (.A1(net2260),
    .A2(net268),
    .B1(net331),
    .B2(net270),
    .C1(_1641_),
    .X(_1642_));
 sky130_fd_sc_hd__mux2_2 _3891_ (.A0(net2301),
    .A1(_1642_),
    .S(net364),
    .X(_1643_));
 sky130_fd_sc_hd__inv_2 _3892_ (.A(_1643_),
    .Y(_1644_));
 sky130_fd_sc_hd__or2_1 _3893_ (.A(_1640_),
    .B(_1643_),
    .X(_1645_));
 sky130_fd_sc_hd__nand2_1 _3894_ (.A(net2377),
    .B(_1643_),
    .Y(_1646_));
 sky130_fd_sc_hd__and2_1 _3895_ (.A(_1645_),
    .B(_1646_),
    .X(_1647_));
 sky130_fd_sc_hd__or4_1 _3896_ (.A(_1611_),
    .B(_1624_),
    .C(_1635_),
    .D(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__or4_2 _3897_ (.A(_1503_),
    .B(_1552_),
    .C(_1600_),
    .D(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__and2b_1 _3898_ (.A_N(net426),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[3] ),
    .X(_1650_));
 sky130_fd_sc_hd__a221o_2 _3899_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[3] ),
    .A2(net361),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[3] ),
    .C1(_1650_),
    .X(_1651_));
 sky130_fd_sc_hd__mux2_2 _3900_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[3] ),
    .A1(_1651_),
    .S(net363),
    .X(_1652_));
 sky130_fd_sc_hd__or2_1 _3901_ (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[3] ),
    .B(net272),
    .X(_1653_));
 sky130_fd_sc_hd__o221a_4 _3902_ (.A1(net610),
    .A2(net274),
    .B1(net244),
    .B2(net330),
    .C1(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__and2_1 _3903_ (.A(net610),
    .B(net346),
    .X(_1655_));
 sky130_fd_sc_hd__a221oi_4 _3904_ (.A1(net2192),
    .A2(net268),
    .B1(net330),
    .B2(net270),
    .C1(_1655_),
    .Y(_1656_));
 sky130_fd_sc_hd__nand2_1 _3905_ (.A(net366),
    .B(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ),
    .Y(_1657_));
 sky130_fd_sc_hd__o21a_1 _3906_ (.A1(net366),
    .A2(_1656_),
    .B1(_1657_),
    .X(_1658_));
 sky130_fd_sc_hd__o21ai_2 _3907_ (.A1(net366),
    .A2(_1656_),
    .B1(_1657_),
    .Y(_1659_));
 sky130_fd_sc_hd__nand2_1 _3908_ (.A(_1654_),
    .B(net201),
    .Y(_1660_));
 sky130_fd_sc_hd__or2_1 _3909_ (.A(_1654_),
    .B(net201),
    .X(_1661_));
 sky130_fd_sc_hd__nand2_1 _3910_ (.A(_1660_),
    .B(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hd__and2b_1 _3911_ (.A_N(net426),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[2] ),
    .X(_1663_));
 sky130_fd_sc_hd__a221o_2 _3912_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[2] ),
    .A2(net361),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[2] ),
    .C1(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__mux2_2 _3913_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[2] ),
    .A1(_1664_),
    .S(net363),
    .X(_1665_));
 sky130_fd_sc_hd__or2_1 _3914_ (.A(net2379),
    .B(net272),
    .X(_1666_));
 sky130_fd_sc_hd__o221a_4 _3915_ (.A1(net923),
    .A2(_1421_),
    .B1(net244),
    .B2(net329),
    .C1(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__and2_1 _3916_ (.A(net923),
    .B(net346),
    .X(_1668_));
 sky130_fd_sc_hd__a221oi_4 _3917_ (.A1(net2160),
    .A2(net268),
    .B1(net329),
    .B2(net270),
    .C1(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hd__nand2_1 _3918_ (.A(net367),
    .B(net2162),
    .Y(_1670_));
 sky130_fd_sc_hd__o21a_1 _3919_ (.A1(net367),
    .A2(_1669_),
    .B1(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__o21ai_1 _3920_ (.A1(net367),
    .A2(_1669_),
    .B1(_1670_),
    .Y(_1672_));
 sky130_fd_sc_hd__xnor2_1 _3921_ (.A(_1667_),
    .B(net197),
    .Y(_1673_));
 sky130_fd_sc_hd__nand2_1 _3922_ (.A(_1662_),
    .B(_1673_),
    .Y(_1674_));
 sky130_fd_sc_hd__and3_1 _3923_ (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(net426),
    .C(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[0] ),
    .X(_1675_));
 sky130_fd_sc_hd__a221o_2 _3924_ (.A1(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[0] ),
    .A2(_1429_),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[0] ),
    .C1(_1675_),
    .X(_1676_));
 sky130_fd_sc_hd__and2_1 _3925_ (.A(net1410),
    .B(net347),
    .X(_1677_));
 sky130_fd_sc_hd__a221oi_4 _3926_ (.A1(net2327),
    .A2(net268),
    .B1(net356),
    .B2(net270),
    .C1(_1677_),
    .Y(_1678_));
 sky130_fd_sc_hd__nand2_1 _3927_ (.A(net367),
    .B(net953),
    .Y(_1679_));
 sky130_fd_sc_hd__o21a_2 _3928_ (.A1(net367),
    .A2(_1678_),
    .B1(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__o21ai_4 _3929_ (.A1(net367),
    .A2(_1678_),
    .B1(_1679_),
    .Y(_1681_));
 sky130_fd_sc_hd__or2_1 _3930_ (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ),
    .B(net272),
    .X(_1682_));
 sky130_fd_sc_hd__o221a_2 _3931_ (.A1(net1410),
    .A2(net274),
    .B1(net244),
    .B2(net356),
    .C1(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__inv_2 _3932_ (.A(_1683_),
    .Y(_1684_));
 sky130_fd_sc_hd__nand2_1 _3933_ (.A(net191),
    .B(_1683_),
    .Y(_1685_));
 sky130_fd_sc_hd__or2_1 _3934_ (.A(net191),
    .B(_1683_),
    .X(_1686_));
 sky130_fd_sc_hd__and2_1 _3935_ (.A(_1685_),
    .B(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__and3_1 _3936_ (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ),
    .B(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .C(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[1] ),
    .X(_1688_));
 sky130_fd_sc_hd__a221o_4 _3937_ (.A1(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[1] ),
    .A2(_1429_),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[1] ),
    .C1(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__inv_2 _3938_ (.A(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__and3b_1 _3939_ (.A_N(net346),
    .B(_1456_),
    .C(_1689_),
    .X(_1691_));
 sky130_fd_sc_hd__and2_1 _3940_ (.A(net1996),
    .B(net347),
    .X(_1692_));
 sky130_fd_sc_hd__and3b_1 _3941_ (.A_N(net346),
    .B(_1457_),
    .C(net2306),
    .X(_1693_));
 sky130_fd_sc_hd__o31a_1 _3942_ (.A1(_1691_),
    .A2(_1692_),
    .A3(_1693_),
    .B1(net364),
    .X(_1694_));
 sky130_fd_sc_hd__nand2_1 _3943_ (.A(net367),
    .B(\U_DATAPATH.U_EX_MEM.i_pc_target_EX[1] ),
    .Y(_1695_));
 sky130_fd_sc_hd__inv_2 _3944_ (.A(_1695_),
    .Y(_1696_));
 sky130_fd_sc_hd__nor2_1 _3945_ (.A(_1694_),
    .B(_1696_),
    .Y(_1697_));
 sky130_fd_sc_hd__or2_1 _3946_ (.A(_1694_),
    .B(_1696_),
    .X(_1698_));
 sky130_fd_sc_hd__or2_1 _3947_ (.A(net2394),
    .B(net272),
    .X(_1699_));
 sky130_fd_sc_hd__o221a_4 _3948_ (.A1(net1996),
    .A2(net274),
    .B1(net244),
    .B2(_1689_),
    .C1(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__inv_2 _3949_ (.A(_1700_),
    .Y(_1701_));
 sky130_fd_sc_hd__or2_1 _3950_ (.A(net186),
    .B(_1700_),
    .X(_1702_));
 sky130_fd_sc_hd__nand2_1 _3951_ (.A(net186),
    .B(_1700_),
    .Y(_1703_));
 sky130_fd_sc_hd__and2b_1 _3952_ (.A_N(net426),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[6] ),
    .X(_1704_));
 sky130_fd_sc_hd__a221o_2 _3953_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[6] ),
    .A2(net361),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[6] ),
    .C1(_1704_),
    .X(_1705_));
 sky130_fd_sc_hd__mux2_1 _3954_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[6] ),
    .A1(_1705_),
    .S(net363),
    .X(_1706_));
 sky130_fd_sc_hd__or2_1 _3955_ (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ),
    .B(net272),
    .X(_1707_));
 sky130_fd_sc_hd__o221a_4 _3956_ (.A1(net1558),
    .A2(net274),
    .B1(net244),
    .B2(net328),
    .C1(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__and2_1 _3957_ (.A(net1558),
    .B(net346),
    .X(_1709_));
 sky130_fd_sc_hd__a221o_2 _3958_ (.A1(net2299),
    .A2(net268),
    .B1(_1706_),
    .B2(net270),
    .C1(_1709_),
    .X(_1710_));
 sky130_fd_sc_hd__mux2_2 _3959_ (.A0(net2244),
    .A1(_1710_),
    .S(net365),
    .X(_1711_));
 sky130_fd_sc_hd__or2_1 _3960_ (.A(_1708_),
    .B(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__nand2_1 _3961_ (.A(_1708_),
    .B(_1711_),
    .Y(_1713_));
 sky130_fd_sc_hd__and2_1 _3962_ (.A(_1712_),
    .B(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__and2b_1 _3963_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[4] ),
    .X(_1715_));
 sky130_fd_sc_hd__a221o_1 _3964_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[4] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[4] ),
    .C1(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__mux2_2 _3965_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[4] ),
    .A1(_1716_),
    .S(net362),
    .X(_1717_));
 sky130_fd_sc_hd__and2_1 _3966_ (.A(net2173),
    .B(net347),
    .X(_1718_));
 sky130_fd_sc_hd__a221o_4 _3967_ (.A1(net2297),
    .A2(net267),
    .B1(net327),
    .B2(net269),
    .C1(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__and2_1 _3968_ (.A(net366),
    .B(net2314),
    .X(_1720_));
 sky130_fd_sc_hd__a21oi_4 _3969_ (.A1(net364),
    .A2(_1719_),
    .B1(_1720_),
    .Y(_1721_));
 sky130_fd_sc_hd__a21o_1 _3970_ (.A1(net364),
    .A2(_1719_),
    .B1(_1720_),
    .X(_1722_));
 sky130_fd_sc_hd__or2_1 _3971_ (.A(net2396),
    .B(net272),
    .X(_1723_));
 sky130_fd_sc_hd__o221a_4 _3972_ (.A1(net2173),
    .A2(net274),
    .B1(net244),
    .B2(_1717_),
    .C1(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__or2_1 _3973_ (.A(net182),
    .B(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__nand2_1 _3974_ (.A(net181),
    .B(_1724_),
    .Y(_1726_));
 sky130_fd_sc_hd__and2b_1 _3975_ (.A_N(net426),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[7] ),
    .X(_1727_));
 sky130_fd_sc_hd__a221o_1 _3976_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[7] ),
    .A2(net361),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[7] ),
    .C1(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__mux2_2 _3977_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[7] ),
    .A1(_1728_),
    .S(net362),
    .X(_1729_));
 sky130_fd_sc_hd__or2_1 _3978_ (.A(net2380),
    .B(net271),
    .X(_1730_));
 sky130_fd_sc_hd__o221a_4 _3979_ (.A1(net1017),
    .A2(net274),
    .B1(net244),
    .B2(_1729_),
    .C1(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__and2_1 _3980_ (.A(net1017),
    .B(net345),
    .X(_1732_));
 sky130_fd_sc_hd__a221o_2 _3981_ (.A1(net2221),
    .A2(net268),
    .B1(net326),
    .B2(net270),
    .C1(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__mux2_2 _3982_ (.A0(net2294),
    .A1(_1733_),
    .S(net364),
    .X(_1734_));
 sky130_fd_sc_hd__or2_1 _3983_ (.A(_1731_),
    .B(_1734_),
    .X(_1735_));
 sky130_fd_sc_hd__nand2_1 _3984_ (.A(_1731_),
    .B(_1734_),
    .Y(_1736_));
 sky130_fd_sc_hd__and2_1 _3985_ (.A(_1735_),
    .B(_1736_),
    .X(_1737_));
 sky130_fd_sc_hd__and2b_1 _3986_ (.A_N(net426),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[5] ),
    .X(_1738_));
 sky130_fd_sc_hd__a221o_4 _3987_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[5] ),
    .A2(net361),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[5] ),
    .C1(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__mux2_1 _3988_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[5] ),
    .A1(_1739_),
    .S(net363),
    .X(_1740_));
 sky130_fd_sc_hd__or2_1 _3989_ (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[5] ),
    .B(net272),
    .X(_1741_));
 sky130_fd_sc_hd__o221a_4 _3990_ (.A1(net660),
    .A2(net274),
    .B1(net244),
    .B2(net325),
    .C1(_1741_),
    .X(_1742_));
 sky130_fd_sc_hd__and2_1 _3991_ (.A(net660),
    .B(net346),
    .X(_1743_));
 sky130_fd_sc_hd__a221o_2 _3992_ (.A1(net2324),
    .A2(net268),
    .B1(net325),
    .B2(net270),
    .C1(_1743_),
    .X(_1744_));
 sky130_fd_sc_hd__mux2_2 _3993_ (.A0(net2388),
    .A1(_1744_),
    .S(net365),
    .X(_1745_));
 sky130_fd_sc_hd__or2_1 _3994_ (.A(_1742_),
    .B(_1745_),
    .X(_1746_));
 sky130_fd_sc_hd__nand2_1 _3995_ (.A(_1742_),
    .B(_1745_),
    .Y(_1747_));
 sky130_fd_sc_hd__and2_1 _3996_ (.A(_1746_),
    .B(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__a2111o_1 _3997_ (.A1(_1725_),
    .A2(_1726_),
    .B1(_1737_),
    .C1(_1748_),
    .D1(_1714_),
    .X(_1749_));
 sky130_fd_sc_hd__and2b_1 _3998_ (.A_N(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[10] ),
    .X(_1750_));
 sky130_fd_sc_hd__a221o_1 _3999_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[10] ),
    .A2(net361),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[10] ),
    .C1(_1750_),
    .X(_1751_));
 sky130_fd_sc_hd__mux2_1 _4000_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[10] ),
    .A1(_1751_),
    .S(net363),
    .X(_1752_));
 sky130_fd_sc_hd__or2_1 _4001_ (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[10] ),
    .B(net272),
    .X(_1753_));
 sky130_fd_sc_hd__o221a_4 _4002_ (.A1(net2033),
    .A2(net274),
    .B1(net244),
    .B2(net324),
    .C1(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__and2_1 _4003_ (.A(net2033),
    .B(net346),
    .X(_1755_));
 sky130_fd_sc_hd__a221o_2 _4004_ (.A1(net2256),
    .A2(net268),
    .B1(_1752_),
    .B2(net270),
    .C1(_1755_),
    .X(_1756_));
 sky130_fd_sc_hd__mux2_2 _4005_ (.A0(net2286),
    .A1(_1756_),
    .S(net365),
    .X(_1757_));
 sky130_fd_sc_hd__or2_1 _4006_ (.A(_1754_),
    .B(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__nand2_1 _4007_ (.A(_1754_),
    .B(_1757_),
    .Y(_1759_));
 sky130_fd_sc_hd__and2_1 _4008_ (.A(_1758_),
    .B(_1759_),
    .X(_1760_));
 sky130_fd_sc_hd__and2b_1 _4009_ (.A_N(net426),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[8] ),
    .X(_1761_));
 sky130_fd_sc_hd__a221o_1 _4010_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[8] ),
    .A2(net361),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[8] ),
    .C1(_1761_),
    .X(_1762_));
 sky130_fd_sc_hd__mux2_2 _4011_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[8] ),
    .A1(_1762_),
    .S(net363),
    .X(_1763_));
 sky130_fd_sc_hd__a22o_1 _4012_ (.A1(net2295),
    .A2(net268),
    .B1(net323),
    .B2(net270),
    .X(_1764_));
 sky130_fd_sc_hd__a21oi_2 _4013_ (.A1(net2133),
    .A2(net347),
    .B1(_1764_),
    .Y(_1765_));
 sky130_fd_sc_hd__nand2_1 _4014_ (.A(net367),
    .B(net2344),
    .Y(_1766_));
 sky130_fd_sc_hd__o21a_1 _4015_ (.A1(net367),
    .A2(_1765_),
    .B1(_1766_),
    .X(_1767_));
 sky130_fd_sc_hd__o21ai_1 _4016_ (.A1(net367),
    .A2(_1765_),
    .B1(_1766_),
    .Y(_1768_));
 sky130_fd_sc_hd__or2_1 _4017_ (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[8] ),
    .B(net272),
    .X(_1769_));
 sky130_fd_sc_hd__o221a_4 _4018_ (.A1(net2133),
    .A2(net274),
    .B1(net244),
    .B2(_1763_),
    .C1(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__or2_1 _4019_ (.A(_1768_),
    .B(_1770_),
    .X(_1771_));
 sky130_fd_sc_hd__nand2_1 _4020_ (.A(_1768_),
    .B(_1770_),
    .Y(_1772_));
 sky130_fd_sc_hd__and2_1 _4021_ (.A(_1771_),
    .B(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__and2b_1 _4022_ (.A_N(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[11] ),
    .X(_1774_));
 sky130_fd_sc_hd__a221o_2 _4023_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[11] ),
    .A2(net361),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[11] ),
    .C1(_1774_),
    .X(_1775_));
 sky130_fd_sc_hd__mux2_1 _4024_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[11] ),
    .A1(_1775_),
    .S(net363),
    .X(_1776_));
 sky130_fd_sc_hd__or2_1 _4025_ (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ),
    .B(net271),
    .X(_1777_));
 sky130_fd_sc_hd__o221a_4 _4026_ (.A1(net2071),
    .A2(net273),
    .B1(net243),
    .B2(_1776_),
    .C1(_1777_),
    .X(_1778_));
 sky130_fd_sc_hd__and2_1 _4027_ (.A(net2071),
    .B(net345),
    .X(_1779_));
 sky130_fd_sc_hd__a221o_2 _4028_ (.A1(net2267),
    .A2(net267),
    .B1(net322),
    .B2(net269),
    .C1(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__mux2_2 _4029_ (.A0(net2397),
    .A1(_1780_),
    .S(net365),
    .X(_1781_));
 sky130_fd_sc_hd__or2_1 _4030_ (.A(_1778_),
    .B(_1781_),
    .X(_1782_));
 sky130_fd_sc_hd__nand2_1 _4031_ (.A(_1778_),
    .B(_1781_),
    .Y(_1783_));
 sky130_fd_sc_hd__and2_1 _4032_ (.A(_1782_),
    .B(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__and2b_1 _4033_ (.A_N(net426),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[9] ),
    .X(_1785_));
 sky130_fd_sc_hd__a221o_1 _4034_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[9] ),
    .A2(net361),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[9] ),
    .C1(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__mux2_2 _4035_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[9] ),
    .A1(_1786_),
    .S(net363),
    .X(_1787_));
 sky130_fd_sc_hd__or2_1 _4036_ (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ),
    .B(net272),
    .X(_1788_));
 sky130_fd_sc_hd__o221a_4 _4037_ (.A1(net2191),
    .A2(_1421_),
    .B1(_1428_),
    .B2(net321),
    .C1(_1788_),
    .X(_1789_));
 sky130_fd_sc_hd__and2_1 _4038_ (.A(net2191),
    .B(net346),
    .X(_1790_));
 sky130_fd_sc_hd__a221o_2 _4039_ (.A1(net2236),
    .A2(net268),
    .B1(_1787_),
    .B2(net270),
    .C1(_1790_),
    .X(_1791_));
 sky130_fd_sc_hd__mux2_2 _4040_ (.A0(net2356),
    .A1(_1791_),
    .S(net365),
    .X(_1792_));
 sky130_fd_sc_hd__inv_2 _4041_ (.A(_1792_),
    .Y(_1793_));
 sky130_fd_sc_hd__or2_1 _4042_ (.A(_1789_),
    .B(_1792_),
    .X(_1794_));
 sky130_fd_sc_hd__nand2_1 _4043_ (.A(_1789_),
    .B(_1792_),
    .Y(_1795_));
 sky130_fd_sc_hd__and2_1 _4044_ (.A(_1794_),
    .B(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__or4_1 _4045_ (.A(_1760_),
    .B(_1773_),
    .C(_1784_),
    .D(_1796_),
    .X(_1797_));
 sky130_fd_sc_hd__and2b_1 _4046_ (.A_N(net426),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[14] ),
    .X(_1798_));
 sky130_fd_sc_hd__a221o_4 _4047_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[14] ),
    .A2(net361),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[14] ),
    .C1(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__mux2_1 _4048_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[14] ),
    .A1(_1799_),
    .S(net363),
    .X(_1800_));
 sky130_fd_sc_hd__or2_1 _4049_ (.A(net2372),
    .B(net272),
    .X(_1801_));
 sky130_fd_sc_hd__o221a_4 _4050_ (.A1(net2066),
    .A2(net274),
    .B1(net244),
    .B2(_1800_),
    .C1(_1801_),
    .X(_1802_));
 sky130_fd_sc_hd__and2_1 _4051_ (.A(net2066),
    .B(net346),
    .X(_1803_));
 sky130_fd_sc_hd__a221o_2 _4052_ (.A1(net2158),
    .A2(net268),
    .B1(net320),
    .B2(net270),
    .C1(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__mux2_2 _4053_ (.A0(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ),
    .A1(_1804_),
    .S(net365),
    .X(_1805_));
 sky130_fd_sc_hd__xor2_1 _4054_ (.A(_1802_),
    .B(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__and2b_1 _4055_ (.A_N(net426),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[12] ),
    .X(_1807_));
 sky130_fd_sc_hd__a221o_1 _4056_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[12] ),
    .A2(net361),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[12] ),
    .C1(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__mux2_2 _4057_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[12] ),
    .A1(_1808_),
    .S(net363),
    .X(_1809_));
 sky130_fd_sc_hd__and2_1 _4058_ (.A(net2137),
    .B(net346),
    .X(_1810_));
 sky130_fd_sc_hd__a221o_1 _4059_ (.A1(net2274),
    .A2(net268),
    .B1(net319),
    .B2(net270),
    .C1(_1810_),
    .X(_1811_));
 sky130_fd_sc_hd__mux2_2 _4060_ (.A0(net2332),
    .A1(_1811_),
    .S(net365),
    .X(_1812_));
 sky130_fd_sc_hd__inv_2 _4061_ (.A(_1812_),
    .Y(_1813_));
 sky130_fd_sc_hd__or2_1 _4062_ (.A(net2369),
    .B(net272),
    .X(_1814_));
 sky130_fd_sc_hd__o221a_4 _4063_ (.A1(net2137),
    .A2(net274),
    .B1(net244),
    .B2(_1809_),
    .C1(_1814_),
    .X(_1815_));
 sky130_fd_sc_hd__or2_1 _4064_ (.A(_1812_),
    .B(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__nand2_1 _4065_ (.A(_1812_),
    .B(net2370),
    .Y(_1817_));
 sky130_fd_sc_hd__and2_1 _4066_ (.A(_1816_),
    .B(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__and2b_1 _4067_ (.A_N(net425),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[15] ),
    .X(_1819_));
 sky130_fd_sc_hd__a221o_2 _4068_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[15] ),
    .A2(net360),
    .B1(net358),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[15] ),
    .C1(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__mux2_1 _4069_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[15] ),
    .A1(_1820_),
    .S(net362),
    .X(_1821_));
 sky130_fd_sc_hd__or2_1 _4070_ (.A(net2384),
    .B(net271),
    .X(_1822_));
 sky130_fd_sc_hd__o221a_4 _4071_ (.A1(net2174),
    .A2(net273),
    .B1(net243),
    .B2(_1821_),
    .C1(_1822_),
    .X(_1823_));
 sky130_fd_sc_hd__and2_1 _4072_ (.A(net2174),
    .B(net345),
    .X(_1824_));
 sky130_fd_sc_hd__a221o_2 _4073_ (.A1(net2302),
    .A2(net267),
    .B1(net318),
    .B2(net269),
    .C1(_1824_),
    .X(_1825_));
 sky130_fd_sc_hd__mux2_2 _4074_ (.A0(net2290),
    .A1(_1825_),
    .S(net364),
    .X(_1826_));
 sky130_fd_sc_hd__or2_1 _4075_ (.A(_1823_),
    .B(_1826_),
    .X(_1827_));
 sky130_fd_sc_hd__nand2_1 _4076_ (.A(net2385),
    .B(_1826_),
    .Y(_1828_));
 sky130_fd_sc_hd__and2_1 _4077_ (.A(_1827_),
    .B(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__and2b_1 _4078_ (.A_N(net426),
    .B(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[13] ),
    .X(_1830_));
 sky130_fd_sc_hd__a221o_1 _4079_ (.A1(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[13] ),
    .A2(net361),
    .B1(net359),
    .B2(\U_DATAPATH.U_MEM_WB.o_read_data_WB[13] ),
    .C1(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__mux2_2 _4080_ (.A0(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[13] ),
    .A1(_1831_),
    .S(net363),
    .X(_1832_));
 sky130_fd_sc_hd__or2_1 _4081_ (.A(net2381),
    .B(net272),
    .X(_1833_));
 sky130_fd_sc_hd__o221a_4 _4082_ (.A1(net1970),
    .A2(net274),
    .B1(net244),
    .B2(net317),
    .C1(_1833_),
    .X(_1834_));
 sky130_fd_sc_hd__and2_1 _4083_ (.A(net1970),
    .B(net346),
    .X(_1835_));
 sky130_fd_sc_hd__a221o_2 _4084_ (.A1(net2240),
    .A2(net268),
    .B1(net317),
    .B2(net270),
    .C1(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__mux2_2 _4085_ (.A0(net2247),
    .A1(_1836_),
    .S(net365),
    .X(_1837_));
 sky130_fd_sc_hd__inv_2 _4086_ (.A(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__or2_1 _4087_ (.A(_1834_),
    .B(_1837_),
    .X(_1839_));
 sky130_fd_sc_hd__nand2_1 _4088_ (.A(_1834_),
    .B(_1837_),
    .Y(_1840_));
 sky130_fd_sc_hd__and2_1 _4089_ (.A(_1839_),
    .B(_1840_),
    .X(_1841_));
 sky130_fd_sc_hd__or4_2 _4090_ (.A(_1806_),
    .B(_1818_),
    .C(_1829_),
    .D(_1841_),
    .X(_1842_));
 sky130_fd_sc_hd__a2111o_1 _4091_ (.A1(_1702_),
    .A2(_1703_),
    .B1(_1797_),
    .C1(_1687_),
    .D1(_1674_),
    .X(_1843_));
 sky130_fd_sc_hd__or4_2 _4092_ (.A(_1649_),
    .B(_1749_),
    .C(_1842_),
    .D(_1843_),
    .X(_1844_));
 sky130_fd_sc_hd__a21oi_1 _4093_ (.A1(net193),
    .A2(_1683_),
    .B1(net189),
    .Y(_1845_));
 sky130_fd_sc_hd__or3_2 _4094_ (.A(net191),
    .B(_1684_),
    .C(net186),
    .X(_1846_));
 sky130_fd_sc_hd__inv_2 _4095_ (.A(_1846_),
    .Y(_1847_));
 sky130_fd_sc_hd__o2111ai_1 _4096_ (.A1(_1701_),
    .A2(_1845_),
    .B1(_1846_),
    .C1(_1673_),
    .D1(_1662_),
    .Y(_1848_));
 sky130_fd_sc_hd__nand2_1 _4097_ (.A(_1662_),
    .B(net196),
    .Y(_1849_));
 sky130_fd_sc_hd__o221a_1 _4098_ (.A1(_1654_),
    .A2(net206),
    .B1(_1667_),
    .B2(_1849_),
    .C1(_1848_),
    .X(_1850_));
 sky130_fd_sc_hd__nand2b_1 _4099_ (.A_N(_1731_),
    .B(_1734_),
    .Y(_1851_));
 sky130_fd_sc_hd__nand2b_1 _4100_ (.A_N(_1708_),
    .B(_1711_),
    .Y(_1852_));
 sky130_fd_sc_hd__nand2b_1 _4101_ (.A_N(_1742_),
    .B(_1745_),
    .Y(_1853_));
 sky130_fd_sc_hd__o31a_1 _4102_ (.A1(net184),
    .A2(_1724_),
    .A3(_1748_),
    .B1(_1853_),
    .X(_1854_));
 sky130_fd_sc_hd__o21a_1 _4103_ (.A1(_1714_),
    .A2(_1854_),
    .B1(_1852_),
    .X(_1855_));
 sky130_fd_sc_hd__o22a_1 _4104_ (.A1(_1749_),
    .A2(_1850_),
    .B1(_1855_),
    .B2(_1737_),
    .X(_1856_));
 sky130_fd_sc_hd__a21o_1 _4105_ (.A1(_1851_),
    .A2(_1856_),
    .B1(_1797_),
    .X(_1857_));
 sky130_fd_sc_hd__nand2b_1 _4106_ (.A_N(_1754_),
    .B(_1757_),
    .Y(_1858_));
 sky130_fd_sc_hd__o32a_1 _4107_ (.A1(_1767_),
    .A2(_1770_),
    .A3(_1796_),
    .B1(_1793_),
    .B2(_1789_),
    .X(_1859_));
 sky130_fd_sc_hd__o21a_1 _4108_ (.A1(_1760_),
    .A2(_1859_),
    .B1(_1858_),
    .X(_1860_));
 sky130_fd_sc_hd__or2_1 _4109_ (.A(_1784_),
    .B(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__nand2b_1 _4110_ (.A_N(_1778_),
    .B(_1781_),
    .Y(_1862_));
 sky130_fd_sc_hd__a31o_1 _4111_ (.A1(_1857_),
    .A2(_1861_),
    .A3(_1862_),
    .B1(_1842_),
    .X(_1863_));
 sky130_fd_sc_hd__nand2b_1 _4112_ (.A_N(_1802_),
    .B(_1805_),
    .Y(_1864_));
 sky130_fd_sc_hd__o32a_1 _4113_ (.A1(_1813_),
    .A2(_1815_),
    .A3(_1841_),
    .B1(_1838_),
    .B2(_1834_),
    .X(_1865_));
 sky130_fd_sc_hd__o21a_1 _4114_ (.A1(_1806_),
    .A2(_1865_),
    .B1(_1864_),
    .X(_1866_));
 sky130_fd_sc_hd__or2_1 _4115_ (.A(_1829_),
    .B(_1866_),
    .X(_1867_));
 sky130_fd_sc_hd__nand2b_1 _4116_ (.A_N(_1823_),
    .B(_1826_),
    .Y(_1868_));
 sky130_fd_sc_hd__a31oi_2 _4117_ (.A1(_1863_),
    .A2(_1867_),
    .A3(_1868_),
    .B1(_1649_),
    .Y(_1869_));
 sky130_fd_sc_hd__nand2_1 _4118_ (.A(_1592_),
    .B(_1595_),
    .Y(_1870_));
 sky130_fd_sc_hd__nand2b_1 _4119_ (.A_N(_1557_),
    .B(_1560_),
    .Y(_1871_));
 sky130_fd_sc_hd__o32a_1 _4120_ (.A1(_1570_),
    .A2(_1572_),
    .A3(_1588_),
    .B1(_1585_),
    .B2(_1580_),
    .X(_1872_));
 sky130_fd_sc_hd__o21a_1 _4121_ (.A1(_1563_),
    .A2(_1872_),
    .B1(_1871_),
    .X(_1873_));
 sky130_fd_sc_hd__nand2b_1 _4122_ (.A_N(_1545_),
    .B(_1548_),
    .Y(_1874_));
 sky130_fd_sc_hd__nand2b_1 _4123_ (.A_N(_1533_),
    .B(_1536_),
    .Y(_1875_));
 sky130_fd_sc_hd__and2b_1 _4124_ (.A_N(_1521_),
    .B(_1526_),
    .X(_1876_));
 sky130_fd_sc_hd__a211oi_1 _4125_ (.A1(_1509_),
    .A2(_1510_),
    .B1(_1513_),
    .C1(_1528_),
    .Y(_1877_));
 sky130_fd_sc_hd__o21ai_1 _4126_ (.A1(_1876_),
    .A2(_1877_),
    .B1(_1539_),
    .Y(_1878_));
 sky130_fd_sc_hd__a21o_1 _4127_ (.A1(_1875_),
    .A2(_1878_),
    .B1(_1551_),
    .X(_1879_));
 sky130_fd_sc_hd__a21o_1 _4128_ (.A1(_1874_),
    .A2(_1879_),
    .B1(_1648_),
    .X(_1880_));
 sky130_fd_sc_hd__nand2b_1 _4129_ (.A_N(_1605_),
    .B(_1608_),
    .Y(_1881_));
 sky130_fd_sc_hd__o32a_1 _4130_ (.A1(_1618_),
    .A2(_1621_),
    .A3(_1647_),
    .B1(_1644_),
    .B2(_1640_),
    .X(_1882_));
 sky130_fd_sc_hd__o21a_1 _4131_ (.A1(_1611_),
    .A2(_1882_),
    .B1(_1881_),
    .X(_1883_));
 sky130_fd_sc_hd__or2_1 _4132_ (.A(_1635_),
    .B(_1883_),
    .X(_1884_));
 sky130_fd_sc_hd__nand2b_1 _4133_ (.A_N(_1629_),
    .B(_1632_),
    .Y(_1885_));
 sky130_fd_sc_hd__a31o_1 _4134_ (.A1(_1880_),
    .A2(_1884_),
    .A3(_1885_),
    .B1(_1503_),
    .X(_1886_));
 sky130_fd_sc_hd__nand2b_1 _4135_ (.A_N(_1471_),
    .B(_1474_),
    .Y(_1887_));
 sky130_fd_sc_hd__o32a_1 _4136_ (.A1(_1466_),
    .A2(_1485_),
    .A3(_1487_),
    .B1(_1463_),
    .B2(_1438_),
    .X(_1888_));
 sky130_fd_sc_hd__o21a_1 _4137_ (.A1(_1477_),
    .A2(_1888_),
    .B1(_1887_),
    .X(_1889_));
 sky130_fd_sc_hd__or2_1 _4138_ (.A(_1501_),
    .B(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__nand2b_1 _4139_ (.A_N(_1494_),
    .B(_1498_),
    .Y(_1891_));
 sky130_fd_sc_hd__a31o_1 _4140_ (.A1(_1886_),
    .A2(_1890_),
    .A3(_1891_),
    .B1(_1600_),
    .X(_1892_));
 sky130_fd_sc_hd__o211ai_2 _4141_ (.A1(_1599_),
    .A2(_1873_),
    .B1(_1892_),
    .C1(_1870_),
    .Y(_1893_));
 sky130_fd_sc_hd__o21ai_2 _4142_ (.A1(_1869_),
    .A2(_1893_),
    .B1(_1844_),
    .Y(_1894_));
 sky130_fd_sc_hd__and3b_1 _4143_ (.A_N(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ),
    .C(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .X(_1895_));
 sky130_fd_sc_hd__xnor2_1 _4144_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .B(_1894_),
    .Y(_1896_));
 sky130_fd_sc_hd__nand3b_2 _4145_ (.A_N(net2340),
    .B(net2315),
    .C(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .Y(_1897_));
 sky130_fd_sc_hd__nand2b_2 _4146_ (.A_N(net2336),
    .B(net2358),
    .Y(_1898_));
 sky130_fd_sc_hd__nand2b_2 _4147_ (.A_N(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .B(net2336),
    .Y(_1899_));
 sky130_fd_sc_hd__or2_2 _4148_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .B(net2315),
    .X(_1900_));
 sky130_fd_sc_hd__o32a_1 _4149_ (.A1(net2340),
    .A2(_1899_),
    .A3(_1900_),
    .B1(_1897_),
    .B2(_1898_),
    .X(_1901_));
 sky130_fd_sc_hd__or3b_2 _4150_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .B(net2340),
    .C_N(net2319),
    .X(_1902_));
 sky130_fd_sc_hd__o21a_1 _4151_ (.A1(_1899_),
    .A2(_1902_),
    .B1(_1901_),
    .X(_1903_));
 sky130_fd_sc_hd__nor2_1 _4152_ (.A(_1844_),
    .B(_1903_),
    .Y(_1904_));
 sky130_fd_sc_hd__nor2_1 _4153_ (.A(_1897_),
    .B(_1899_),
    .Y(_1905_));
 sky130_fd_sc_hd__a221o_1 _4154_ (.A1(_1895_),
    .A2(_1896_),
    .B1(_1905_),
    .B2(_1844_),
    .C1(_1904_),
    .X(_1906_));
 sky130_fd_sc_hd__a21oi_1 _4155_ (.A1(net2248),
    .A2(_1906_),
    .B1(net2114),
    .Y(_1907_));
 sky130_fd_sc_hd__xor2_1 _4156_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ),
    .B(net2203),
    .X(_1908_));
 sky130_fd_sc_hd__a21oi_1 _4157_ (.A1(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ),
    .A2(net2130),
    .B1(_1908_),
    .Y(_1909_));
 sky130_fd_sc_hd__and3_1 _4158_ (.A(net2162),
    .B(net2130),
    .C(_1908_),
    .X(_1910_));
 sky130_fd_sc_hd__nor2_1 _4159_ (.A(net2131),
    .B(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__mux2_2 _4160_ (.A0(net2132),
    .A1(net2024),
    .S(net176),
    .X(_1912_));
 sky130_fd_sc_hd__xor2_1 _4161_ (.A(net2162),
    .B(net2130),
    .X(_1913_));
 sky130_fd_sc_hd__mux2_2 _4162_ (.A0(_1913_),
    .A1(net2122),
    .S(net179),
    .X(_1914_));
 sky130_fd_sc_hd__inv_2 _4163_ (.A(_1914_),
    .Y(_1915_));
 sky130_fd_sc_hd__nand2_1 _4164_ (.A(_1912_),
    .B(_1914_),
    .Y(_1916_));
 sky130_fd_sc_hd__a21oi_1 _4165_ (.A1(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ),
    .A2(net2203),
    .B1(_1910_),
    .Y(_1917_));
 sky130_fd_sc_hd__nor2_1 _4166_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ),
    .B(\U_DATAPATH.U_ID_EX.o_pc_EX[4] ),
    .Y(_1918_));
 sky130_fd_sc_hd__nand2_1 _4167_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ),
    .B(\U_DATAPATH.U_ID_EX.o_pc_EX[4] ),
    .Y(_1919_));
 sky130_fd_sc_hd__and2b_1 _4168_ (.A_N(_1918_),
    .B(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__xnor2_1 _4169_ (.A(net2204),
    .B(_1920_),
    .Y(_1921_));
 sky130_fd_sc_hd__mux2_1 _4170_ (.A0(net2205),
    .A1(net2068),
    .S(net173),
    .X(_1922_));
 sky130_fd_sc_hd__nand2b_1 _4171_ (.A_N(_1916_),
    .B(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hd__or2_1 _4172_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ),
    .B(net2206),
    .X(_1924_));
 sky130_fd_sc_hd__nand2_1 _4173_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ),
    .B(net2206),
    .Y(_1925_));
 sky130_fd_sc_hd__nand2_1 _4174_ (.A(_1924_),
    .B(net2207),
    .Y(_1926_));
 sky130_fd_sc_hd__o21a_1 _4175_ (.A1(net2204),
    .A2(_1918_),
    .B1(_1919_),
    .X(_1927_));
 sky130_fd_sc_hd__xor2_1 _4176_ (.A(net2208),
    .B(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__mux2_1 _4177_ (.A0(net2209),
    .A1(net837),
    .S(net176),
    .X(_1929_));
 sky130_fd_sc_hd__nand2b_2 _4178_ (.A_N(_1923_),
    .B(_1929_),
    .Y(_1930_));
 sky130_fd_sc_hd__o21a_1 _4179_ (.A1(_1926_),
    .A2(_1927_),
    .B1(net2207),
    .X(_1931_));
 sky130_fd_sc_hd__nor2_1 _4180_ (.A(net2244),
    .B(net2216),
    .Y(_1932_));
 sky130_fd_sc_hd__nand2_1 _4181_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ),
    .B(net2216),
    .Y(_1933_));
 sky130_fd_sc_hd__and2b_1 _4182_ (.A_N(_1932_),
    .B(net2217),
    .X(_1934_));
 sky130_fd_sc_hd__xnor2_1 _4183_ (.A(_1931_),
    .B(_1934_),
    .Y(_1935_));
 sky130_fd_sc_hd__mux2_1 _4184_ (.A0(_1935_),
    .A1(net817),
    .S(net176),
    .X(_1936_));
 sky130_fd_sc_hd__inv_2 _4185_ (.A(_1936_),
    .Y(_1937_));
 sky130_fd_sc_hd__nor2_1 _4186_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ),
    .B(net2140),
    .Y(_1938_));
 sky130_fd_sc_hd__nand2_1 _4187_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ),
    .B(net2140),
    .Y(_1939_));
 sky130_fd_sc_hd__nand2b_1 _4188_ (.A_N(_1938_),
    .B(net2141),
    .Y(_1940_));
 sky130_fd_sc_hd__o21a_1 _4189_ (.A1(_1931_),
    .A2(_1932_),
    .B1(net2217),
    .X(_1941_));
 sky130_fd_sc_hd__xor2_1 _4190_ (.A(_1940_),
    .B(net2218),
    .X(_1942_));
 sky130_fd_sc_hd__mux2_1 _4191_ (.A0(_1942_),
    .A1(net2065),
    .S(net176),
    .X(_1943_));
 sky130_fd_sc_hd__inv_2 _4192_ (.A(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__or3_1 _4193_ (.A(_1930_),
    .B(_1937_),
    .C(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__nor2_1 _4194_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ),
    .B(\U_DATAPATH.U_ID_EX.o_pc_EX[8] ),
    .Y(_1946_));
 sky130_fd_sc_hd__nand2_1 _4195_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ),
    .B(\U_DATAPATH.U_ID_EX.o_pc_EX[8] ),
    .Y(_1947_));
 sky130_fd_sc_hd__nand2b_1 _4196_ (.A_N(_1946_),
    .B(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__o21a_1 _4197_ (.A1(_1938_),
    .A2(_1941_),
    .B1(net2141),
    .X(_1949_));
 sky130_fd_sc_hd__xor2_1 _4198_ (.A(_1948_),
    .B(net2142),
    .X(_1950_));
 sky130_fd_sc_hd__mux2_1 _4199_ (.A0(net2143),
    .A1(net1893),
    .S(net179),
    .X(_1951_));
 sky130_fd_sc_hd__nand2b_1 _4200_ (.A_N(_1945_),
    .B(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__nor2_1 _4201_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ),
    .B(net2231),
    .Y(_1953_));
 sky130_fd_sc_hd__nand2_1 _4202_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ),
    .B(net2231),
    .Y(_1954_));
 sky130_fd_sc_hd__nand2b_1 _4203_ (.A_N(_1953_),
    .B(net2232),
    .Y(_1955_));
 sky130_fd_sc_hd__o21a_1 _4204_ (.A1(_1946_),
    .A2(net2142),
    .B1(_1947_),
    .X(_1956_));
 sky130_fd_sc_hd__xor2_1 _4205_ (.A(net2233),
    .B(_1956_),
    .X(_1957_));
 sky130_fd_sc_hd__mux2_1 _4206_ (.A0(net2234),
    .A1(net1998),
    .S(net178),
    .X(_1958_));
 sky130_fd_sc_hd__nand2b_1 _4207_ (.A_N(_1952_),
    .B(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__nor2_1 _4208_ (.A(net2286),
    .B(net2052),
    .Y(_1960_));
 sky130_fd_sc_hd__nand2_1 _4209_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[10] ),
    .B(net2052),
    .Y(_1961_));
 sky130_fd_sc_hd__nand2b_1 _4210_ (.A_N(_1960_),
    .B(net2053),
    .Y(_1962_));
 sky130_fd_sc_hd__o21a_1 _4211_ (.A1(_1953_),
    .A2(_1956_),
    .B1(net2232),
    .X(_1963_));
 sky130_fd_sc_hd__xor2_1 _4212_ (.A(_1962_),
    .B(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__mux2_1 _4213_ (.A0(_1964_),
    .A1(net1994),
    .S(net178),
    .X(_1965_));
 sky130_fd_sc_hd__and2b_1 _4214_ (.A_N(_1959_),
    .B(_1965_),
    .X(_1966_));
 sky130_fd_sc_hd__nor2_1 _4215_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ),
    .B(net2316),
    .Y(_1967_));
 sky130_fd_sc_hd__nand2_1 _4216_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ),
    .B(net2316),
    .Y(_1968_));
 sky130_fd_sc_hd__nand2b_1 _4217_ (.A_N(_1967_),
    .B(_1968_),
    .Y(_1969_));
 sky130_fd_sc_hd__o21a_1 _4218_ (.A1(_1960_),
    .A2(_1963_),
    .B1(net2053),
    .X(_1970_));
 sky130_fd_sc_hd__xor2_1 _4219_ (.A(_1969_),
    .B(net2054),
    .X(_1971_));
 sky130_fd_sc_hd__mux2_1 _4220_ (.A0(_1971_),
    .A1(net2022),
    .S(net178),
    .X(_1972_));
 sky130_fd_sc_hd__nor2_1 _4221_ (.A(net2332),
    .B(net2184),
    .Y(_1973_));
 sky130_fd_sc_hd__nand2_1 _4222_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ),
    .B(net2184),
    .Y(_1974_));
 sky130_fd_sc_hd__nand2b_1 _4223_ (.A_N(_1973_),
    .B(net2185),
    .Y(_1975_));
 sky130_fd_sc_hd__o21a_1 _4224_ (.A1(_1967_),
    .A2(net2054),
    .B1(net2317),
    .X(_1976_));
 sky130_fd_sc_hd__xor2_1 _4225_ (.A(_1975_),
    .B(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__mux2_1 _4226_ (.A0(_1977_),
    .A1(net2003),
    .S(net178),
    .X(_1978_));
 sky130_fd_sc_hd__and3_1 _4227_ (.A(_1966_),
    .B(_1972_),
    .C(_1978_),
    .X(_1979_));
 sky130_fd_sc_hd__nor2_1 _4228_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ),
    .B(net2163),
    .Y(_1980_));
 sky130_fd_sc_hd__nand2_1 _4229_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ),
    .B(net2163),
    .Y(_1981_));
 sky130_fd_sc_hd__nand2b_1 _4230_ (.A_N(_1980_),
    .B(net2164),
    .Y(_1982_));
 sky130_fd_sc_hd__o21a_1 _4231_ (.A1(_1973_),
    .A2(_1976_),
    .B1(net2185),
    .X(_1983_));
 sky130_fd_sc_hd__xor2_1 _4232_ (.A(_1982_),
    .B(net2186),
    .X(_1984_));
 sky130_fd_sc_hd__mux2_1 _4233_ (.A0(_1984_),
    .A1(net1792),
    .S(net178),
    .X(_1985_));
 sky130_fd_sc_hd__nand2_1 _4234_ (.A(net2005),
    .B(_1985_),
    .Y(_1986_));
 sky130_fd_sc_hd__nor2_1 _4235_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ),
    .B(\U_DATAPATH.U_ID_EX.o_pc_EX[14] ),
    .Y(_1987_));
 sky130_fd_sc_hd__nand2_1 _4236_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ),
    .B(\U_DATAPATH.U_ID_EX.o_pc_EX[14] ),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2b_1 _4237_ (.A_N(_1987_),
    .B(_1988_),
    .Y(_1989_));
 sky130_fd_sc_hd__o21a_1 _4238_ (.A1(_1980_),
    .A2(_1983_),
    .B1(net2164),
    .X(_1990_));
 sky130_fd_sc_hd__xor2_1 _4239_ (.A(_1989_),
    .B(net2165),
    .X(_1991_));
 sky130_fd_sc_hd__mux2_1 _4240_ (.A0(net2166),
    .A1(net1242),
    .S(net178),
    .X(_1992_));
 sky130_fd_sc_hd__and3_4 _4241_ (.A(_1979_),
    .B(_1985_),
    .C(_1992_),
    .X(_1993_));
 sky130_fd_sc_hd__nor2_1 _4242_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ),
    .B(net2060),
    .Y(_1994_));
 sky130_fd_sc_hd__nand2_1 _4243_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ),
    .B(net2060),
    .Y(_1995_));
 sky130_fd_sc_hd__nand2b_1 _4244_ (.A_N(_1994_),
    .B(net2061),
    .Y(_1996_));
 sky130_fd_sc_hd__o21a_2 _4245_ (.A1(_1987_),
    .A2(_1990_),
    .B1(_1988_),
    .X(_1997_));
 sky130_fd_sc_hd__xor2_1 _4246_ (.A(net2062),
    .B(_1997_),
    .X(_1998_));
 sky130_fd_sc_hd__mux2_1 _4247_ (.A0(net2063),
    .A1(net2036),
    .S(net169),
    .X(_1999_));
 sky130_fd_sc_hd__and2_1 _4248_ (.A(_1993_),
    .B(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__nor2_1 _4249_ (.A(net2212),
    .B(\U_DATAPATH.U_ID_EX.o_pc_EX[16] ),
    .Y(_2001_));
 sky130_fd_sc_hd__nand2_1 _4250_ (.A(net2212),
    .B(\U_DATAPATH.U_ID_EX.o_pc_EX[16] ),
    .Y(_2002_));
 sky130_fd_sc_hd__nand2b_1 _4251_ (.A_N(_2001_),
    .B(net2213),
    .Y(_2003_));
 sky130_fd_sc_hd__o21a_1 _4252_ (.A1(_1994_),
    .A2(_1997_),
    .B1(net2061),
    .X(_2004_));
 sky130_fd_sc_hd__xor2_1 _4253_ (.A(net2214),
    .B(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__mux2_1 _4254_ (.A0(_2005_),
    .A1(net1997),
    .S(net169),
    .X(_2006_));
 sky130_fd_sc_hd__nand2_1 _4255_ (.A(_2000_),
    .B(_2006_),
    .Y(_2007_));
 sky130_fd_sc_hd__nor2_1 _4256_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ),
    .B(net2040),
    .Y(_2008_));
 sky130_fd_sc_hd__nand2_1 _4257_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ),
    .B(net2040),
    .Y(_2009_));
 sky130_fd_sc_hd__nand2b_1 _4258_ (.A_N(_2008_),
    .B(net2041),
    .Y(_2010_));
 sky130_fd_sc_hd__o21a_1 _4259_ (.A1(_2001_),
    .A2(_2004_),
    .B1(_2002_),
    .X(_2011_));
 sky130_fd_sc_hd__xor2_1 _4260_ (.A(net2042),
    .B(_2011_),
    .X(_2012_));
 sky130_fd_sc_hd__mux2_1 _4261_ (.A0(net2043),
    .A1(net1984),
    .S(net169),
    .X(_2013_));
 sky130_fd_sc_hd__and3_1 _4262_ (.A(_2000_),
    .B(_2006_),
    .C(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__nor2_1 _4263_ (.A(net2235),
    .B(net2012),
    .Y(_2015_));
 sky130_fd_sc_hd__nand2_1 _4264_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[18] ),
    .B(net2012),
    .Y(_2016_));
 sky130_fd_sc_hd__nand2b_1 _4265_ (.A_N(_2015_),
    .B(net2013),
    .Y(_2017_));
 sky130_fd_sc_hd__o21a_1 _4266_ (.A1(_2008_),
    .A2(_2011_),
    .B1(net2041),
    .X(_2018_));
 sky130_fd_sc_hd__xor2_1 _4267_ (.A(net2014),
    .B(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__mux2_1 _4268_ (.A0(net2015),
    .A1(net1987),
    .S(net171),
    .X(_2020_));
 sky130_fd_sc_hd__and2_1 _4269_ (.A(_2014_),
    .B(_2020_),
    .X(_2021_));
 sky130_fd_sc_hd__nor2_1 _4270_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ),
    .B(net2177),
    .Y(_2022_));
 sky130_fd_sc_hd__nand2_1 _4271_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ),
    .B(net2177),
    .Y(_2023_));
 sky130_fd_sc_hd__nand2b_1 _4272_ (.A_N(_2022_),
    .B(net2178),
    .Y(_2024_));
 sky130_fd_sc_hd__o21a_1 _4273_ (.A1(_2015_),
    .A2(_2018_),
    .B1(net2013),
    .X(_2025_));
 sky130_fd_sc_hd__xor2_1 _4274_ (.A(net2179),
    .B(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__mux2_1 _4275_ (.A0(_2026_),
    .A1(net1784),
    .S(net170),
    .X(_2027_));
 sky130_fd_sc_hd__nand2_1 _4276_ (.A(_2021_),
    .B(_2027_),
    .Y(_2028_));
 sky130_fd_sc_hd__nor2_1 _4277_ (.A(net2325),
    .B(net2320),
    .Y(_2029_));
 sky130_fd_sc_hd__nand2_1 _4278_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ),
    .B(net2320),
    .Y(_2030_));
 sky130_fd_sc_hd__nand2b_1 _4279_ (.A_N(_2029_),
    .B(net2321),
    .Y(_2031_));
 sky130_fd_sc_hd__o21a_1 _4280_ (.A1(_2022_),
    .A2(_2025_),
    .B1(net2178),
    .X(_2032_));
 sky130_fd_sc_hd__xor2_1 _4281_ (.A(_2031_),
    .B(_2032_),
    .X(_2033_));
 sky130_fd_sc_hd__mux2_1 _4282_ (.A0(_2033_),
    .A1(net2019),
    .S(net171),
    .X(_2034_));
 sky130_fd_sc_hd__and3_1 _4283_ (.A(_2021_),
    .B(_2027_),
    .C(_2034_),
    .X(_2035_));
 sky130_fd_sc_hd__nor2_1 _4284_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ),
    .B(net2276),
    .Y(_2036_));
 sky130_fd_sc_hd__nand2_1 _4285_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ),
    .B(net2276),
    .Y(_2037_));
 sky130_fd_sc_hd__nand2b_1 _4286_ (.A_N(_2036_),
    .B(net2277),
    .Y(_2038_));
 sky130_fd_sc_hd__o21a_1 _4287_ (.A1(_2029_),
    .A2(_2032_),
    .B1(_2030_),
    .X(_2039_));
 sky130_fd_sc_hd__xor2_1 _4288_ (.A(net2278),
    .B(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__mux2_1 _4289_ (.A0(net2279),
    .A1(net1969),
    .S(net170),
    .X(_2041_));
 sky130_fd_sc_hd__and2_1 _4290_ (.A(_2035_),
    .B(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__nor2_1 _4291_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ),
    .B(net2227),
    .Y(_2043_));
 sky130_fd_sc_hd__nand2_1 _4292_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ),
    .B(net2227),
    .Y(_2044_));
 sky130_fd_sc_hd__nand2b_1 _4293_ (.A_N(_2043_),
    .B(net2228),
    .Y(_2045_));
 sky130_fd_sc_hd__o21a_1 _4294_ (.A1(_2036_),
    .A2(_2039_),
    .B1(_2037_),
    .X(_2046_));
 sky130_fd_sc_hd__xor2_1 _4295_ (.A(net2229),
    .B(_2046_),
    .X(_2047_));
 sky130_fd_sc_hd__mux2_1 _4296_ (.A0(net2230),
    .A1(net1820),
    .S(net169),
    .X(_2048_));
 sky130_fd_sc_hd__nand2_1 _4297_ (.A(_2042_),
    .B(_2048_),
    .Y(_2049_));
 sky130_fd_sc_hd__nor2_1 _4298_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ),
    .B(net2270),
    .Y(_2050_));
 sky130_fd_sc_hd__nand2_1 _4299_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ),
    .B(net2270),
    .Y(_2051_));
 sky130_fd_sc_hd__nand2b_1 _4300_ (.A_N(_2050_),
    .B(net2271),
    .Y(_2052_));
 sky130_fd_sc_hd__o21a_1 _4301_ (.A1(_2043_),
    .A2(_2046_),
    .B1(net2228),
    .X(_2053_));
 sky130_fd_sc_hd__xnor2_1 _4302_ (.A(net2272),
    .B(_2053_),
    .Y(_2054_));
 sky130_fd_sc_hd__inv_2 _4303_ (.A(net2273),
    .Y(_2055_));
 sky130_fd_sc_hd__mux2_1 _4304_ (.A0(_2055_),
    .A1(net2038),
    .S(net169),
    .X(_2056_));
 sky130_fd_sc_hd__and3_1 _4305_ (.A(_2042_),
    .B(_2048_),
    .C(_2056_),
    .X(_2057_));
 sky130_fd_sc_hd__or2_1 _4306_ (.A(net2151),
    .B(\U_DATAPATH.U_ID_EX.o_pc_EX[24] ),
    .X(_2058_));
 sky130_fd_sc_hd__nand2_1 _4307_ (.A(net2151),
    .B(\U_DATAPATH.U_ID_EX.o_pc_EX[24] ),
    .Y(_2059_));
 sky130_fd_sc_hd__nand2_1 _4308_ (.A(_2058_),
    .B(net2152),
    .Y(_2060_));
 sky130_fd_sc_hd__o21a_1 _4309_ (.A1(_2050_),
    .A2(_2053_),
    .B1(net2271),
    .X(_2061_));
 sky130_fd_sc_hd__xor2_1 _4310_ (.A(net2153),
    .B(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__mux2_1 _4311_ (.A0(net2154),
    .A1(net2000),
    .S(net171),
    .X(_2063_));
 sky130_fd_sc_hd__nand2_1 _4312_ (.A(_2057_),
    .B(_2063_),
    .Y(_2064_));
 sky130_fd_sc_hd__or2_1 _4313_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ),
    .B(net2309),
    .X(_2065_));
 sky130_fd_sc_hd__nand2_1 _4314_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ),
    .B(net2309),
    .Y(_2066_));
 sky130_fd_sc_hd__nand2_1 _4315_ (.A(_2065_),
    .B(net2310),
    .Y(_2067_));
 sky130_fd_sc_hd__o21a_1 _4316_ (.A1(net2153),
    .A2(_2061_),
    .B1(net2152),
    .X(_2068_));
 sky130_fd_sc_hd__xnor2_1 _4317_ (.A(net2311),
    .B(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__inv_2 _4318_ (.A(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__mux2_1 _4319_ (.A0(_2070_),
    .A1(net2017),
    .S(net171),
    .X(_2071_));
 sky130_fd_sc_hd__and3_1 _4320_ (.A(_2057_),
    .B(_2063_),
    .C(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__o21a_1 _4321_ (.A1(_2067_),
    .A2(_2068_),
    .B1(_2066_),
    .X(_2073_));
 sky130_fd_sc_hd__nor2_1 _4322_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ),
    .B(net2223),
    .Y(_2074_));
 sky130_fd_sc_hd__nand2_1 _4323_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ),
    .B(net2223),
    .Y(_2075_));
 sky130_fd_sc_hd__and2b_1 _4324_ (.A_N(_2074_),
    .B(net2224),
    .X(_2076_));
 sky130_fd_sc_hd__xnor2_1 _4325_ (.A(_2073_),
    .B(net2225),
    .Y(_2077_));
 sky130_fd_sc_hd__mux2_1 _4326_ (.A0(net2226),
    .A1(net1993),
    .S(net171),
    .X(_2078_));
 sky130_fd_sc_hd__and4_2 _4327_ (.A(_2057_),
    .B(_2063_),
    .C(_2071_),
    .D(_2078_),
    .X(_2079_));
 sky130_fd_sc_hd__nor2_1 _4328_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ),
    .B(net2194),
    .Y(_2080_));
 sky130_fd_sc_hd__nand2_1 _4329_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ),
    .B(net2194),
    .Y(_2081_));
 sky130_fd_sc_hd__nand2b_1 _4330_ (.A_N(_2080_),
    .B(net2195),
    .Y(_2082_));
 sky130_fd_sc_hd__o21a_1 _4331_ (.A1(_2073_),
    .A2(_2074_),
    .B1(_2075_),
    .X(_2083_));
 sky130_fd_sc_hd__xor2_1 _4332_ (.A(net2196),
    .B(_2083_),
    .X(_2084_));
 sky130_fd_sc_hd__mux2_2 _4333_ (.A0(net2197),
    .A1(net871),
    .S(net172),
    .X(_2085_));
 sky130_fd_sc_hd__nand2_1 _4334_ (.A(_2079_),
    .B(_2085_),
    .Y(_2086_));
 sky130_fd_sc_hd__nor2_1 _4335_ (.A(net2201),
    .B(net2029),
    .Y(_2087_));
 sky130_fd_sc_hd__nand2_1 _4336_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[28] ),
    .B(net2029),
    .Y(_2088_));
 sky130_fd_sc_hd__nand2b_1 _4337_ (.A_N(_2087_),
    .B(net2030),
    .Y(_2089_));
 sky130_fd_sc_hd__o21a_1 _4338_ (.A1(_2080_),
    .A2(_2083_),
    .B1(net2195),
    .X(_2090_));
 sky130_fd_sc_hd__xor2_1 _4339_ (.A(_2089_),
    .B(_2090_),
    .X(_2091_));
 sky130_fd_sc_hd__mux2_1 _4340_ (.A0(_2091_),
    .A1(net2011),
    .S(net172),
    .X(_2092_));
 sky130_fd_sc_hd__nand3_1 _4341_ (.A(_2079_),
    .B(_2085_),
    .C(_2092_),
    .Y(_2093_));
 sky130_fd_sc_hd__nor2_1 _4342_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ),
    .B(net2249),
    .Y(_2094_));
 sky130_fd_sc_hd__nand2_1 _4343_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ),
    .B(net2249),
    .Y(_2095_));
 sky130_fd_sc_hd__nand2b_1 _4344_ (.A_N(_2094_),
    .B(_2095_),
    .Y(_2096_));
 sky130_fd_sc_hd__o21a_1 _4345_ (.A1(_2087_),
    .A2(_2090_),
    .B1(net2030),
    .X(_2097_));
 sky130_fd_sc_hd__xor2_1 _4346_ (.A(_2096_),
    .B(net2031),
    .X(_2098_));
 sky130_fd_sc_hd__mux2_1 _4347_ (.A0(_2098_),
    .A1(net2008),
    .S(net172),
    .X(_2099_));
 sky130_fd_sc_hd__or2_1 _4348_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ),
    .B(\U_DATAPATH.U_ID_EX.o_pc_EX[30] ),
    .X(_2100_));
 sky130_fd_sc_hd__nand2_1 _4349_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ),
    .B(\U_DATAPATH.U_ID_EX.o_pc_EX[30] ),
    .Y(_2101_));
 sky130_fd_sc_hd__nand2_1 _4350_ (.A(_2100_),
    .B(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__o21a_1 _4351_ (.A1(_2094_),
    .A2(net2031),
    .B1(net2250),
    .X(_2103_));
 sky130_fd_sc_hd__xor2_1 _4352_ (.A(_2102_),
    .B(net2251),
    .X(_2104_));
 sky130_fd_sc_hd__mux2_1 _4353_ (.A0(net2252),
    .A1(net1983),
    .S(net172),
    .X(_2105_));
 sky130_fd_sc_hd__and3b_1 _4354_ (.A_N(_2093_),
    .B(_2099_),
    .C(_2105_),
    .X(_2106_));
 sky130_fd_sc_hd__o21a_1 _4355_ (.A1(_2102_),
    .A2(_2103_),
    .B1(_2101_),
    .X(_2107_));
 sky130_fd_sc_hd__xor2_1 _4356_ (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ),
    .B(net2025),
    .X(_2108_));
 sky130_fd_sc_hd__xnor2_1 _4357_ (.A(_2107_),
    .B(net2026),
    .Y(_2109_));
 sky130_fd_sc_hd__mux2_1 _4358_ (.A0(net2027),
    .A1(net1990),
    .S(net173),
    .X(_2110_));
 sky130_fd_sc_hd__xnor2_1 _4359_ (.A(net385),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .Y(_2111_));
 sky130_fd_sc_hd__a2bb2o_1 _4360_ (.A1_N(_1402_),
    .A2_N(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .B1(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .B2(_1400_),
    .X(_2112_));
 sky130_fd_sc_hd__a221o_1 _4361_ (.A1(_1402_),
    .A2(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .B1(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .B2(_1401_),
    .C1(_2112_),
    .X(_2113_));
 sky130_fd_sc_hd__o221ai_1 _4362_ (.A1(_1401_),
    .A2(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .B1(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .B2(_1400_),
    .C1(_2111_),
    .Y(_2114_));
 sky130_fd_sc_hd__xor2_1 _4363_ (.A(net424),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .X(_2115_));
 sky130_fd_sc_hd__xor2_1 _4364_ (.A(net399),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .X(_2116_));
 sky130_fd_sc_hd__xor2_1 _4365_ (.A(net414),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .X(_2117_));
 sky130_fd_sc_hd__xor2_1 _4366_ (.A(net404),
    .B(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .X(_2118_));
 sky130_fd_sc_hd__or4_1 _4367_ (.A(_2115_),
    .B(_2116_),
    .C(_2117_),
    .D(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__o21a_1 _4368_ (.A1(_2113_),
    .A2(_2114_),
    .B1(_2119_),
    .X(_2120_));
 sky130_fd_sc_hd__nor3b_1 _4369_ (.A(net1716),
    .B(_2120_),
    .C_N(net1342),
    .Y(_2121_));
 sky130_fd_sc_hd__or3b_1 _4370_ (.A(net1716),
    .B(_2120_),
    .C_N(net1342),
    .X(_2122_));
 sky130_fd_sc_hd__nor2_1 _4371_ (.A(_2106_),
    .B(net236),
    .Y(_2123_));
 sky130_fd_sc_hd__nand2_1 _4372_ (.A(_2106_),
    .B(net2028),
    .Y(_2124_));
 sky130_fd_sc_hd__o21a_1 _4373_ (.A1(_2106_),
    .A2(_2110_),
    .B1(net222),
    .X(_2125_));
 sky130_fd_sc_hd__a22o_1 _4374_ (.A1(net1990),
    .A2(net237),
    .B1(_2124_),
    .B2(_2125_),
    .X(_1267_));
 sky130_fd_sc_hd__a41o_1 _4375_ (.A1(_2079_),
    .A2(_2085_),
    .A3(_2092_),
    .A4(_2099_),
    .B1(_2105_),
    .X(_2126_));
 sky130_fd_sc_hd__a22o_1 _4376_ (.A1(net1983),
    .A2(net236),
    .B1(_2123_),
    .B2(_2126_),
    .X(_1266_));
 sky130_fd_sc_hd__xnor2_1 _4377_ (.A(_2093_),
    .B(_2099_),
    .Y(_2127_));
 sky130_fd_sc_hd__mux2_1 _4378_ (.A0(net2008),
    .A1(_2127_),
    .S(net220),
    .X(_1265_));
 sky130_fd_sc_hd__and2_1 _4379_ (.A(net2011),
    .B(net236),
    .X(_2128_));
 sky130_fd_sc_hd__a21o_1 _4380_ (.A1(_2079_),
    .A2(_2085_),
    .B1(_2092_),
    .X(_2129_));
 sky130_fd_sc_hd__a31o_1 _4381_ (.A1(_2093_),
    .A2(net220),
    .A3(_2129_),
    .B1(_2128_),
    .X(_1264_));
 sky130_fd_sc_hd__and2_1 _4382_ (.A(net871),
    .B(net236),
    .X(_2130_));
 sky130_fd_sc_hd__or2_1 _4383_ (.A(_2079_),
    .B(_2085_),
    .X(_2131_));
 sky130_fd_sc_hd__a31o_1 _4384_ (.A1(_2086_),
    .A2(net220),
    .A3(_2131_),
    .B1(_2130_),
    .X(_1263_));
 sky130_fd_sc_hd__xor2_1 _4385_ (.A(_2072_),
    .B(_2078_),
    .X(_2132_));
 sky130_fd_sc_hd__mux2_1 _4386_ (.A0(net1993),
    .A1(_2132_),
    .S(net219),
    .X(_1262_));
 sky130_fd_sc_hd__xnor2_1 _4387_ (.A(_2064_),
    .B(net2018),
    .Y(_2133_));
 sky130_fd_sc_hd__mux2_1 _4388_ (.A0(net2017),
    .A1(_2133_),
    .S(net218),
    .X(_1261_));
 sky130_fd_sc_hd__and2_1 _4389_ (.A(net2000),
    .B(net235),
    .X(_2134_));
 sky130_fd_sc_hd__or2_1 _4390_ (.A(_2057_),
    .B(_2063_),
    .X(_2135_));
 sky130_fd_sc_hd__a31o_1 _4391_ (.A1(_2064_),
    .A2(net218),
    .A3(_2135_),
    .B1(_2134_),
    .X(_1260_));
 sky130_fd_sc_hd__xnor2_1 _4392_ (.A(_2049_),
    .B(_2056_),
    .Y(_2136_));
 sky130_fd_sc_hd__mux2_1 _4393_ (.A0(net2038),
    .A1(_2136_),
    .S(net214),
    .X(_1259_));
 sky130_fd_sc_hd__and2_1 _4394_ (.A(net1820),
    .B(net233),
    .X(_2137_));
 sky130_fd_sc_hd__or2_1 _4395_ (.A(_2042_),
    .B(_2048_),
    .X(_2138_));
 sky130_fd_sc_hd__a31o_1 _4396_ (.A1(_2049_),
    .A2(net215),
    .A3(_2138_),
    .B1(_2137_),
    .X(_1258_));
 sky130_fd_sc_hd__or2_1 _4397_ (.A(_2035_),
    .B(_2041_),
    .X(_2139_));
 sky130_fd_sc_hd__nor2_1 _4398_ (.A(_2042_),
    .B(net234),
    .Y(_2140_));
 sky130_fd_sc_hd__a22o_1 _4399_ (.A1(net1969),
    .A2(net234),
    .B1(net2021),
    .B2(_2140_),
    .X(_1257_));
 sky130_fd_sc_hd__a31o_1 _4400_ (.A1(_2014_),
    .A2(_2020_),
    .A3(_2027_),
    .B1(net2020),
    .X(_2141_));
 sky130_fd_sc_hd__nor2_1 _4401_ (.A(_2035_),
    .B(net234),
    .Y(_2142_));
 sky130_fd_sc_hd__a22o_1 _4402_ (.A1(net2019),
    .A2(net237),
    .B1(_2141_),
    .B2(_2142_),
    .X(_1256_));
 sky130_fd_sc_hd__and2_1 _4403_ (.A(net1784),
    .B(net234),
    .X(_2143_));
 sky130_fd_sc_hd__or2_1 _4404_ (.A(_2021_),
    .B(_2027_),
    .X(_2144_));
 sky130_fd_sc_hd__a31o_1 _4405_ (.A1(_2028_),
    .A2(net219),
    .A3(_2144_),
    .B1(_2143_),
    .X(_1255_));
 sky130_fd_sc_hd__or2_1 _4406_ (.A(_2014_),
    .B(_2020_),
    .X(_2145_));
 sky130_fd_sc_hd__nor2_1 _4407_ (.A(_2021_),
    .B(net234),
    .Y(_2146_));
 sky130_fd_sc_hd__a22o_1 _4408_ (.A1(net1987),
    .A2(net235),
    .B1(_2145_),
    .B2(_2146_),
    .X(_1254_));
 sky130_fd_sc_hd__a31o_1 _4409_ (.A1(_1993_),
    .A2(_1999_),
    .A3(_2006_),
    .B1(_2013_),
    .X(_2147_));
 sky130_fd_sc_hd__nor2_1 _4410_ (.A(_2014_),
    .B(net233),
    .Y(_2148_));
 sky130_fd_sc_hd__a22o_1 _4411_ (.A1(net1984),
    .A2(net233),
    .B1(_2147_),
    .B2(_2148_),
    .X(_1253_));
 sky130_fd_sc_hd__and2_1 _4412_ (.A(net1997),
    .B(net233),
    .X(_2149_));
 sky130_fd_sc_hd__or2_1 _4413_ (.A(_2000_),
    .B(_2006_),
    .X(_2150_));
 sky130_fd_sc_hd__a31o_1 _4414_ (.A1(_2007_),
    .A2(net214),
    .A3(_2150_),
    .B1(_2149_),
    .X(_1252_));
 sky130_fd_sc_hd__or2_1 _4415_ (.A(_1993_),
    .B(_1999_),
    .X(_2151_));
 sky130_fd_sc_hd__nor2_1 _4416_ (.A(_2000_),
    .B(net233),
    .Y(_2152_));
 sky130_fd_sc_hd__a22o_1 _4417_ (.A1(net2036),
    .A2(net233),
    .B1(_2151_),
    .B2(_2152_),
    .X(_1251_));
 sky130_fd_sc_hd__a21o_1 _4418_ (.A1(net2005),
    .A2(_1985_),
    .B1(_1992_),
    .X(_2153_));
 sky130_fd_sc_hd__nor2_1 _4419_ (.A(_1993_),
    .B(net240),
    .Y(_2154_));
 sky130_fd_sc_hd__a22o_1 _4420_ (.A1(net1242),
    .A2(net240),
    .B1(net2006),
    .B2(_2154_),
    .X(_1250_));
 sky130_fd_sc_hd__and2_1 _4421_ (.A(net1792),
    .B(net240),
    .X(_2155_));
 sky130_fd_sc_hd__or2_1 _4422_ (.A(_1979_),
    .B(_1985_),
    .X(_2156_));
 sky130_fd_sc_hd__a31o_1 _4423_ (.A1(_1986_),
    .A2(net230),
    .A3(_2156_),
    .B1(_2155_),
    .X(_1249_));
 sky130_fd_sc_hd__a21o_1 _4424_ (.A1(_1966_),
    .A2(net2056),
    .B1(net2004),
    .X(_2157_));
 sky130_fd_sc_hd__nor2_1 _4425_ (.A(net2005),
    .B(net240),
    .Y(_2158_));
 sky130_fd_sc_hd__a22o_1 _4426_ (.A1(net2003),
    .A2(net240),
    .B1(_2157_),
    .B2(_2158_),
    .X(_1248_));
 sky130_fd_sc_hd__or2_1 _4427_ (.A(_1966_),
    .B(net2056),
    .X(_2159_));
 sky130_fd_sc_hd__a21oi_1 _4428_ (.A1(_1966_),
    .A2(net2056),
    .B1(net240),
    .Y(_2160_));
 sky130_fd_sc_hd__a22o_1 _4429_ (.A1(net2022),
    .A2(net241),
    .B1(_2159_),
    .B2(_2160_),
    .X(_1247_));
 sky130_fd_sc_hd__xnor2_1 _4430_ (.A(_1959_),
    .B(_1965_),
    .Y(_2161_));
 sky130_fd_sc_hd__mux2_1 _4431_ (.A0(net1994),
    .A1(_2161_),
    .S(net231),
    .X(_1246_));
 sky130_fd_sc_hd__xnor2_1 _4432_ (.A(_1952_),
    .B(_1958_),
    .Y(_2162_));
 sky130_fd_sc_hd__mux2_1 _4433_ (.A0(net1998),
    .A1(_2162_),
    .S(net230),
    .X(_1245_));
 sky130_fd_sc_hd__and2_1 _4434_ (.A(net1893),
    .B(net238),
    .X(_2163_));
 sky130_fd_sc_hd__nand2b_1 _4435_ (.A_N(_1951_),
    .B(_1945_),
    .Y(_2164_));
 sky130_fd_sc_hd__a31o_1 _4436_ (.A1(_1952_),
    .A2(net227),
    .A3(_2164_),
    .B1(_2163_),
    .X(_1244_));
 sky130_fd_sc_hd__and2_1 _4437_ (.A(net2065),
    .B(net238),
    .X(_2165_));
 sky130_fd_sc_hd__o21ai_1 _4438_ (.A1(_1930_),
    .A2(_1937_),
    .B1(_1944_),
    .Y(_2166_));
 sky130_fd_sc_hd__a31o_1 _4439_ (.A1(_1945_),
    .A2(net226),
    .A3(_2166_),
    .B1(_2165_),
    .X(_1243_));
 sky130_fd_sc_hd__xnor2_1 _4440_ (.A(_1930_),
    .B(_1936_),
    .Y(_2167_));
 sky130_fd_sc_hd__mux2_1 _4441_ (.A0(net817),
    .A1(_2167_),
    .S(net226),
    .X(_1242_));
 sky130_fd_sc_hd__and2_1 _4442_ (.A(net837),
    .B(net238),
    .X(_2168_));
 sky130_fd_sc_hd__a31o_1 _4443_ (.A1(_1912_),
    .A2(_1914_),
    .A3(_1922_),
    .B1(_1929_),
    .X(_2169_));
 sky130_fd_sc_hd__a31o_1 _4444_ (.A1(_1930_),
    .A2(net226),
    .A3(_2169_),
    .B1(_2168_),
    .X(_1241_));
 sky130_fd_sc_hd__and2_1 _4445_ (.A(net2068),
    .B(net236),
    .X(_2170_));
 sky130_fd_sc_hd__a21o_1 _4446_ (.A1(_1912_),
    .A2(_1914_),
    .B1(_1922_),
    .X(_2171_));
 sky130_fd_sc_hd__a31o_1 _4447_ (.A1(_1923_),
    .A2(net221),
    .A3(_2171_),
    .B1(_2170_),
    .X(_1240_));
 sky130_fd_sc_hd__and2_1 _4448_ (.A(net2024),
    .B(net238),
    .X(_2172_));
 sky130_fd_sc_hd__or2_1 _4449_ (.A(_1912_),
    .B(_1914_),
    .X(_2173_));
 sky130_fd_sc_hd__a31o_1 _4450_ (.A1(_1916_),
    .A2(net226),
    .A3(_2173_),
    .B1(_2172_),
    .X(_1239_));
 sky130_fd_sc_hd__mux2_1 _4451_ (.A0(net2122),
    .A1(_1915_),
    .S(net226),
    .X(_1238_));
 sky130_fd_sc_hd__and2_1 _4452_ (.A(\U_DATAPATH.U_EX_MEM.o_mem_write_M ),
    .B(net427),
    .X(_1043_));
 sky130_fd_sc_hd__and2_1 _4453_ (.A(net435),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[31] ),
    .X(_1042_));
 sky130_fd_sc_hd__and2_1 _4454_ (.A(net451),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[30] ),
    .X(_1041_));
 sky130_fd_sc_hd__and2_1 _4455_ (.A(net429),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[29] ),
    .X(_1040_));
 sky130_fd_sc_hd__and2_1 _4456_ (.A(net428),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[28] ),
    .X(_1039_));
 sky130_fd_sc_hd__and2_1 _4457_ (.A(net427),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[27] ),
    .X(_1038_));
 sky130_fd_sc_hd__and2_1 _4458_ (.A(net427),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[26] ),
    .X(_1037_));
 sky130_fd_sc_hd__and2_1 _4459_ (.A(net439),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[25] ),
    .X(_1036_));
 sky130_fd_sc_hd__and2_1 _4460_ (.A(net457),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[24] ),
    .X(_1035_));
 sky130_fd_sc_hd__and2_1 _4461_ (.A(net435),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[23] ),
    .X(_1034_));
 sky130_fd_sc_hd__and2_1 _4462_ (.A(net454),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[22] ),
    .X(_1033_));
 sky130_fd_sc_hd__and2_1 _4463_ (.A(net428),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[21] ),
    .X(_1032_));
 sky130_fd_sc_hd__and2_1 _4464_ (.A(net427),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[20] ),
    .X(_1031_));
 sky130_fd_sc_hd__and2_1 _4465_ (.A(net432),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[19] ),
    .X(_1030_));
 sky130_fd_sc_hd__and2_1 _4466_ (.A(net454),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[18] ),
    .X(_1029_));
 sky130_fd_sc_hd__and2_1 _4467_ (.A(net449),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[17] ),
    .X(_1028_));
 sky130_fd_sc_hd__and2_1 _4468_ (.A(net433),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[16] ),
    .X(_1027_));
 sky130_fd_sc_hd__and2_1 _4469_ (.A(net427),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[15] ),
    .X(_1026_));
 sky130_fd_sc_hd__and2_1 _4470_ (.A(net427),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[14] ),
    .X(_1025_));
 sky130_fd_sc_hd__and2_1 _4471_ (.A(net428),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[13] ),
    .X(_1024_));
 sky130_fd_sc_hd__and2_1 _4472_ (.A(net448),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[12] ),
    .X(_1023_));
 sky130_fd_sc_hd__and2_1 _4473_ (.A(net445),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[11] ),
    .X(_1022_));
 sky130_fd_sc_hd__and2_1 _4474_ (.A(net457),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[10] ),
    .X(_1021_));
 sky130_fd_sc_hd__and2_1 _4475_ (.A(net448),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[9] ),
    .X(_1020_));
 sky130_fd_sc_hd__and2_1 _4476_ (.A(net445),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[8] ),
    .X(_1019_));
 sky130_fd_sc_hd__and2_1 _4477_ (.A(net436),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[7] ),
    .X(_1018_));
 sky130_fd_sc_hd__and2_1 _4478_ (.A(net447),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[6] ),
    .X(_1017_));
 sky130_fd_sc_hd__and2_1 _4479_ (.A(net447),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[5] ),
    .X(_1016_));
 sky130_fd_sc_hd__and2_1 _4480_ (.A(net454),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[4] ),
    .X(_1015_));
 sky130_fd_sc_hd__and2_1 _4481_ (.A(net432),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[3] ),
    .X(_1014_));
 sky130_fd_sc_hd__and2_1 _4482_ (.A(net435),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[2] ),
    .X(_1013_));
 sky130_fd_sc_hd__and2_1 _4483_ (.A(net433),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[1] ),
    .X(_1012_));
 sky130_fd_sc_hd__and2_1 _4484_ (.A(net438),
    .B(\U_DATAPATH.U_EX_MEM.o_write_data_M[0] ),
    .X(_1011_));
 sky130_fd_sc_hd__mux2_1 _4485_ (.A0(net2098),
    .A1(net2028),
    .S(net222),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _4486_ (.A0(net2070),
    .A1(_2105_),
    .S(net222),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _4487_ (.A0(net2093),
    .A1(net2009),
    .S(net220),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _4488_ (.A0(net2096),
    .A1(_2092_),
    .S(net220),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _4489_ (.A0(net2097),
    .A1(_2085_),
    .S(net220),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _4490_ (.A0(net2080),
    .A1(_2078_),
    .S(net217),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _4491_ (.A0(net2082),
    .A1(net2018),
    .S(net218),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _4492_ (.A0(net2067),
    .A1(_2063_),
    .S(net218),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _4493_ (.A0(net2069),
    .A1(_2056_),
    .S(net214),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _4494_ (.A0(net2034),
    .A1(_2048_),
    .S(net215),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _4495_ (.A0(net2047),
    .A1(_2041_),
    .S(net217),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _4496_ (.A0(net2059),
    .A1(net2020),
    .S(net218),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _4497_ (.A0(net2078),
    .A1(_2027_),
    .S(net220),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _4498_ (.A0(net2075),
    .A1(_2020_),
    .S(net216),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _4499_ (.A0(net2086),
    .A1(_2013_),
    .S(net214),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _4500_ (.A0(net2089),
    .A1(_2006_),
    .S(net214),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _4501_ (.A0(net2108),
    .A1(_1999_),
    .S(net214),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _4502_ (.A0(net2088),
    .A1(_1992_),
    .S(net231),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _4503_ (.A0(net2046),
    .A1(_1985_),
    .S(net230),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _4504_ (.A0(net2079),
    .A1(net2004),
    .S(net231),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _4505_ (.A0(net2081),
    .A1(net2023),
    .S(net228),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _4506_ (.A0(net2074),
    .A1(_1965_),
    .S(net227),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _4507_ (.A0(net2073),
    .A1(_1958_),
    .S(net230),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _4508_ (.A0(net2064),
    .A1(net2144),
    .S(net227),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _4509_ (.A0(net2044),
    .A1(net2220),
    .S(net225),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _4510_ (.A0(net2103),
    .A1(_1936_),
    .S(net226),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _4511_ (.A0(net2058),
    .A1(_1929_),
    .S(net226),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _4512_ (.A0(net2072),
    .A1(_1922_),
    .S(net221),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _4513_ (.A0(net2051),
    .A1(_1912_),
    .S(net226),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _4514_ (.A0(net2057),
    .A1(_1914_),
    .S(net225),
    .X(_0292_));
 sky130_fd_sc_hd__nand2b_4 _4515_ (.A_N(net2210),
    .B(net2254),
    .Y(_2174_));
 sky130_fd_sc_hd__and3b_1 _4516_ (.A_N(net2258),
    .B(net2170),
    .C(net1988),
    .X(_2175_));
 sky130_fd_sc_hd__nand2b_2 _4517_ (.A_N(_2174_),
    .B(_2175_),
    .Y(_2176_));
 sky130_fd_sc_hd__or3b_4 _4518_ (.A(net1988),
    .B(net2170),
    .C_N(net2258),
    .X(_2177_));
 sky130_fd_sc_hd__o21a_1 _4519_ (.A1(_2174_),
    .A2(_2177_),
    .B1(_2176_),
    .X(_3636_));
 sky130_fd_sc_hd__mux4_1 _4520_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ),
    .S0(net396),
    .S1(net385),
    .X(_2178_));
 sky130_fd_sc_hd__mux4_1 _4521_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ),
    .S0(net396),
    .S1(net385),
    .X(_2179_));
 sky130_fd_sc_hd__mux2_1 _4522_ (.A0(_2178_),
    .A1(_2179_),
    .S(net375),
    .X(_2180_));
 sky130_fd_sc_hd__mux4_1 _4523_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ),
    .S1(net385),
    .X(_2181_));
 sky130_fd_sc_hd__mux4_1 _4524_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ),
    .S0(net396),
    .S1(net385),
    .X(_2182_));
 sky130_fd_sc_hd__mux2_1 _4525_ (.A0(_2182_),
    .A1(_2181_),
    .S(net375),
    .X(_2183_));
 sky130_fd_sc_hd__mux2_1 _4526_ (.A0(_2183_),
    .A1(_2180_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .X(_0000_));
 sky130_fd_sc_hd__mux4_1 _4527_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ),
    .S0(net396),
    .S1(net385),
    .X(_2184_));
 sky130_fd_sc_hd__mux4_1 _4528_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ),
    .S0(net396),
    .S1(net385),
    .X(_2185_));
 sky130_fd_sc_hd__mux2_1 _4529_ (.A0(_2184_),
    .A1(_2185_),
    .S(net375),
    .X(_2186_));
 sky130_fd_sc_hd__mux4_1 _4530_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ),
    .S0(net396),
    .S1(net385),
    .X(_2187_));
 sky130_fd_sc_hd__mux4_1 _4531_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ),
    .S1(net385),
    .X(_2188_));
 sky130_fd_sc_hd__mux2_1 _4532_ (.A0(_2188_),
    .A1(_2187_),
    .S(net375),
    .X(_2189_));
 sky130_fd_sc_hd__mux2_1 _4533_ (.A0(_2189_),
    .A1(_2186_),
    .S(net369),
    .X(_0011_));
 sky130_fd_sc_hd__mux4_1 _4534_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ),
    .S0(net395),
    .S1(net383),
    .X(_2190_));
 sky130_fd_sc_hd__mux4_1 _4535_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ),
    .S0(net395),
    .S1(net383),
    .X(_2191_));
 sky130_fd_sc_hd__mux2_1 _4536_ (.A0(_2190_),
    .A1(_2191_),
    .S(net374),
    .X(_2192_));
 sky130_fd_sc_hd__mux4_1 _4537_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ),
    .S0(net396),
    .S1(net385),
    .X(_2193_));
 sky130_fd_sc_hd__mux4_1 _4538_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ),
    .S0(net395),
    .S1(net385),
    .X(_2194_));
 sky130_fd_sc_hd__mux2_1 _4539_ (.A0(_2194_),
    .A1(_2193_),
    .S(net375),
    .X(_2195_));
 sky130_fd_sc_hd__mux2_1 _4540_ (.A0(_2195_),
    .A1(_2192_),
    .S(net369),
    .X(_0022_));
 sky130_fd_sc_hd__mux4_1 _4541_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ),
    .S0(net395),
    .S1(net382),
    .X(_2196_));
 sky130_fd_sc_hd__mux4_1 _4542_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ),
    .S0(net395),
    .S1(net383),
    .X(_2197_));
 sky130_fd_sc_hd__mux2_1 _4543_ (.A0(_2196_),
    .A1(_2197_),
    .S(net374),
    .X(_2198_));
 sky130_fd_sc_hd__mux4_1 _4544_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ),
    .S0(net394),
    .S1(net382),
    .X(_2199_));
 sky130_fd_sc_hd__mux4_1 _4545_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ),
    .S0(net394),
    .S1(net383),
    .X(_2200_));
 sky130_fd_sc_hd__mux2_1 _4546_ (.A0(_2200_),
    .A1(_2199_),
    .S(net373),
    .X(_2201_));
 sky130_fd_sc_hd__mux2_1 _4547_ (.A0(_2201_),
    .A1(_2198_),
    .S(net369),
    .X(_0025_));
 sky130_fd_sc_hd__mux4_1 _4548_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ),
    .S0(net391),
    .S1(net380),
    .X(_2202_));
 sky130_fd_sc_hd__mux4_1 _4549_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ),
    .S0(net391),
    .S1(net380),
    .X(_2203_));
 sky130_fd_sc_hd__mux2_1 _4550_ (.A0(_2202_),
    .A1(_2203_),
    .S(net372),
    .X(_2204_));
 sky130_fd_sc_hd__mux4_1 _4551_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ),
    .S0(net391),
    .S1(net380),
    .X(_2205_));
 sky130_fd_sc_hd__mux4_1 _4552_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ),
    .S0(net391),
    .S1(net380),
    .X(_2206_));
 sky130_fd_sc_hd__mux2_1 _4553_ (.A0(_2206_),
    .A1(_2205_),
    .S(net372),
    .X(_2207_));
 sky130_fd_sc_hd__mux2_1 _4554_ (.A0(_2207_),
    .A1(_2204_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .X(_0026_));
 sky130_fd_sc_hd__mux4_1 _4555_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ),
    .S0(net392),
    .S1(net381),
    .X(_2208_));
 sky130_fd_sc_hd__mux4_1 _4556_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ),
    .S0(net392),
    .S1(net381),
    .X(_2209_));
 sky130_fd_sc_hd__mux2_1 _4557_ (.A0(_2208_),
    .A1(_2209_),
    .S(net373),
    .X(_2210_));
 sky130_fd_sc_hd__mux4_1 _4558_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ),
    .S0(net392),
    .S1(net381),
    .X(_2211_));
 sky130_fd_sc_hd__mux4_1 _4559_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ),
    .S0(net392),
    .S1(net381),
    .X(_2212_));
 sky130_fd_sc_hd__mux2_1 _4560_ (.A0(_2212_),
    .A1(_2211_),
    .S(net373),
    .X(_2213_));
 sky130_fd_sc_hd__mux2_1 _4561_ (.A0(_2213_),
    .A1(_2210_),
    .S(net369),
    .X(_0027_));
 sky130_fd_sc_hd__mux4_1 _4562_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ),
    .S0(net394),
    .S1(net382),
    .X(_2214_));
 sky130_fd_sc_hd__mux4_1 _4563_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ),
    .S0(net394),
    .S1(net382),
    .X(_2215_));
 sky130_fd_sc_hd__mux2_1 _4564_ (.A0(_2214_),
    .A1(_2215_),
    .S(net373),
    .X(_2216_));
 sky130_fd_sc_hd__mux4_1 _4565_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ),
    .S0(net394),
    .S1(net382),
    .X(_2217_));
 sky130_fd_sc_hd__mux4_1 _4566_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ),
    .S0(net394),
    .S1(net382),
    .X(_2218_));
 sky130_fd_sc_hd__mux2_1 _4567_ (.A0(_2218_),
    .A1(_2217_),
    .S(net373),
    .X(_2219_));
 sky130_fd_sc_hd__mux2_1 _4568_ (.A0(_2219_),
    .A1(_2216_),
    .S(net369),
    .X(_0028_));
 sky130_fd_sc_hd__mux4_1 _4569_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ),
    .S1(net386),
    .X(_2220_));
 sky130_fd_sc_hd__mux4_1 _4570_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ),
    .S1(net380),
    .X(_2221_));
 sky130_fd_sc_hd__mux2_1 _4571_ (.A0(_2220_),
    .A1(_2221_),
    .S(net372),
    .X(_2222_));
 sky130_fd_sc_hd__mux4_1 _4572_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ),
    .S0(net391),
    .S1(net380),
    .X(_2223_));
 sky130_fd_sc_hd__mux4_1 _4573_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ),
    .S0(net391),
    .S1(net386),
    .X(_2224_));
 sky130_fd_sc_hd__mux2_1 _4574_ (.A0(_2224_),
    .A1(_2223_),
    .S(net372),
    .X(_2225_));
 sky130_fd_sc_hd__mux2_1 _4575_ (.A0(_2225_),
    .A1(_2222_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .X(_0029_));
 sky130_fd_sc_hd__mux4_1 _4576_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ),
    .S0(net396),
    .S1(net385),
    .X(_2226_));
 sky130_fd_sc_hd__mux4_1 _4577_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ),
    .S0(net396),
    .S1(net386),
    .X(_2227_));
 sky130_fd_sc_hd__mux2_1 _4578_ (.A0(_2226_),
    .A1(_2227_),
    .S(net375),
    .X(_2228_));
 sky130_fd_sc_hd__mux4_1 _4579_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ),
    .S0(net396),
    .S1(net385),
    .X(_2229_));
 sky130_fd_sc_hd__mux4_1 _4580_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ),
    .S0(net396),
    .S1(net385),
    .X(_2230_));
 sky130_fd_sc_hd__mux2_1 _4581_ (.A0(_2230_),
    .A1(_2229_),
    .S(net375),
    .X(_2231_));
 sky130_fd_sc_hd__mux2_1 _4582_ (.A0(_2231_),
    .A1(_2228_),
    .S(net369),
    .X(_0030_));
 sky130_fd_sc_hd__mux4_1 _4583_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ),
    .S0(net394),
    .S1(net382),
    .X(_2232_));
 sky130_fd_sc_hd__mux4_1 _4584_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ),
    .S0(net394),
    .S1(net382),
    .X(_2233_));
 sky130_fd_sc_hd__mux2_1 _4585_ (.A0(_2232_),
    .A1(_2233_),
    .S(net374),
    .X(_2234_));
 sky130_fd_sc_hd__mux4_1 _4586_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ),
    .S0(net394),
    .S1(net382),
    .X(_2235_));
 sky130_fd_sc_hd__mux4_1 _4587_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ),
    .S0(net394),
    .S1(net382),
    .X(_2236_));
 sky130_fd_sc_hd__mux2_1 _4588_ (.A0(_2236_),
    .A1(_2235_),
    .S(net374),
    .X(_2237_));
 sky130_fd_sc_hd__mux2_1 _4589_ (.A0(_2237_),
    .A1(_2234_),
    .S(net369),
    .X(_0031_));
 sky130_fd_sc_hd__mux4_1 _4590_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ),
    .S0(net394),
    .S1(net382),
    .X(_2238_));
 sky130_fd_sc_hd__mux4_1 _4591_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ),
    .S0(net394),
    .S1(net382),
    .X(_2239_));
 sky130_fd_sc_hd__mux2_1 _4592_ (.A0(_2238_),
    .A1(_2239_),
    .S(net373),
    .X(_2240_));
 sky130_fd_sc_hd__mux4_1 _4593_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ),
    .S0(net394),
    .S1(net382),
    .X(_2241_));
 sky130_fd_sc_hd__mux4_1 _4594_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ),
    .S0(net394),
    .S1(net382),
    .X(_2242_));
 sky130_fd_sc_hd__mux2_1 _4595_ (.A0(_2242_),
    .A1(_2241_),
    .S(net374),
    .X(_2243_));
 sky130_fd_sc_hd__mux2_1 _4596_ (.A0(_2243_),
    .A1(_2240_),
    .S(net369),
    .X(_0001_));
 sky130_fd_sc_hd__mux4_1 _4597_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ),
    .S0(net389),
    .S1(net378),
    .X(_2244_));
 sky130_fd_sc_hd__mux4_1 _4598_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ),
    .S0(net389),
    .S1(net378),
    .X(_2245_));
 sky130_fd_sc_hd__mux2_1 _4599_ (.A0(_2244_),
    .A1(_2245_),
    .S(net371),
    .X(_2246_));
 sky130_fd_sc_hd__mux4_1 _4600_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ),
    .S0(net389),
    .S1(net378),
    .X(_2247_));
 sky130_fd_sc_hd__mux4_1 _4601_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ),
    .S0(net389),
    .S1(net378),
    .X(_2248_));
 sky130_fd_sc_hd__mux2_1 _4602_ (.A0(_2248_),
    .A1(_2247_),
    .S(net370),
    .X(_2249_));
 sky130_fd_sc_hd__mux2_1 _4603_ (.A0(_2249_),
    .A1(_2246_),
    .S(net368),
    .X(_0002_));
 sky130_fd_sc_hd__mux4_1 _4604_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ),
    .S0(net395),
    .S1(net383),
    .X(_2250_));
 sky130_fd_sc_hd__mux4_1 _4605_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ),
    .S0(net395),
    .S1(net382),
    .X(_2251_));
 sky130_fd_sc_hd__mux2_1 _4606_ (.A0(_2250_),
    .A1(_2251_),
    .S(net374),
    .X(_2252_));
 sky130_fd_sc_hd__mux4_1 _4607_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ),
    .S0(net395),
    .S1(net383),
    .X(_2253_));
 sky130_fd_sc_hd__mux4_1 _4608_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ),
    .S0(net395),
    .S1(net383),
    .X(_2254_));
 sky130_fd_sc_hd__mux2_1 _4609_ (.A0(_2254_),
    .A1(_2253_),
    .S(net374),
    .X(_2255_));
 sky130_fd_sc_hd__mux2_1 _4610_ (.A0(_2255_),
    .A1(_2252_),
    .S(net369),
    .X(_0003_));
 sky130_fd_sc_hd__mux4_1 _4611_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ),
    .S0(net395),
    .S1(net384),
    .X(_2256_));
 sky130_fd_sc_hd__mux4_1 _4612_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ),
    .S0(net393),
    .S1(net384),
    .X(_2257_));
 sky130_fd_sc_hd__mux2_1 _4613_ (.A0(_2256_),
    .A1(_2257_),
    .S(net373),
    .X(_2258_));
 sky130_fd_sc_hd__mux4_1 _4614_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ),
    .S0(net393),
    .S1(net384),
    .X(_2259_));
 sky130_fd_sc_hd__mux4_1 _4615_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ),
    .S0(net393),
    .S1(net384),
    .X(_2260_));
 sky130_fd_sc_hd__mux2_1 _4616_ (.A0(_2260_),
    .A1(_2259_),
    .S(net373),
    .X(_2261_));
 sky130_fd_sc_hd__mux2_1 _4617_ (.A0(_2261_),
    .A1(_2258_),
    .S(net369),
    .X(_0004_));
 sky130_fd_sc_hd__mux4_1 _4618_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ),
    .S0(net392),
    .S1(net381),
    .X(_2262_));
 sky130_fd_sc_hd__mux4_1 _4619_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ),
    .S0(net392),
    .S1(net384),
    .X(_2263_));
 sky130_fd_sc_hd__mux2_1 _4620_ (.A0(_2262_),
    .A1(_2263_),
    .S(net373),
    .X(_2264_));
 sky130_fd_sc_hd__mux4_1 _4621_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ),
    .S0(net392),
    .S1(net381),
    .X(_2265_));
 sky130_fd_sc_hd__mux4_1 _4622_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ),
    .S0(net392),
    .S1(net381),
    .X(_2266_));
 sky130_fd_sc_hd__mux2_1 _4623_ (.A0(_2266_),
    .A1(_2265_),
    .S(net373),
    .X(_2267_));
 sky130_fd_sc_hd__mux2_1 _4624_ (.A0(_2267_),
    .A1(_2264_),
    .S(net369),
    .X(_0005_));
 sky130_fd_sc_hd__mux4_1 _4625_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ),
    .S0(net387),
    .S1(net376),
    .X(_2268_));
 sky130_fd_sc_hd__mux4_1 _4626_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ),
    .S0(net387),
    .S1(net376),
    .X(_2269_));
 sky130_fd_sc_hd__mux2_1 _4627_ (.A0(_2268_),
    .A1(_2269_),
    .S(net370),
    .X(_2270_));
 sky130_fd_sc_hd__mux4_1 _4628_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ),
    .S0(net387),
    .S1(net376),
    .X(_2271_));
 sky130_fd_sc_hd__mux4_1 _4629_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ),
    .S0(net387),
    .S1(net376),
    .X(_2272_));
 sky130_fd_sc_hd__mux2_1 _4630_ (.A0(_2272_),
    .A1(_2271_),
    .S(net370),
    .X(_2273_));
 sky130_fd_sc_hd__mux2_1 _4631_ (.A0(_2273_),
    .A1(_2270_),
    .S(net368),
    .X(_0006_));
 sky130_fd_sc_hd__mux4_1 _4632_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ),
    .S0(net389),
    .S1(net378),
    .X(_2274_));
 sky130_fd_sc_hd__mux4_1 _4633_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ),
    .S0(net392),
    .S1(net381),
    .X(_2275_));
 sky130_fd_sc_hd__mux2_1 _4634_ (.A0(_2274_),
    .A1(_2275_),
    .S(net371),
    .X(_2276_));
 sky130_fd_sc_hd__mux4_1 _4635_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ),
    .S0(net389),
    .S1(net378),
    .X(_2277_));
 sky130_fd_sc_hd__mux4_1 _4636_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ),
    .S0(net389),
    .S1(net378),
    .X(_2278_));
 sky130_fd_sc_hd__mux2_1 _4637_ (.A0(_2278_),
    .A1(_2277_),
    .S(net371),
    .X(_2279_));
 sky130_fd_sc_hd__mux2_1 _4638_ (.A0(_2279_),
    .A1(_2276_),
    .S(net368),
    .X(_0007_));
 sky130_fd_sc_hd__mux4_1 _4639_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ),
    .S0(net394),
    .S1(net382),
    .X(_2280_));
 sky130_fd_sc_hd__mux4_1 _4640_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ),
    .S0(net394),
    .S1(net383),
    .X(_2281_));
 sky130_fd_sc_hd__mux2_1 _4641_ (.A0(_2280_),
    .A1(_2281_),
    .S(net374),
    .X(_2282_));
 sky130_fd_sc_hd__mux4_1 _4642_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ),
    .S0(net392),
    .S1(net381),
    .X(_2283_));
 sky130_fd_sc_hd__mux4_1 _4643_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ),
    .S0(net392),
    .S1(net384),
    .X(_2284_));
 sky130_fd_sc_hd__mux2_1 _4644_ (.A0(_2284_),
    .A1(_2283_),
    .S(net373),
    .X(_2285_));
 sky130_fd_sc_hd__mux2_1 _4645_ (.A0(_2285_),
    .A1(_2282_),
    .S(net369),
    .X(_0008_));
 sky130_fd_sc_hd__mux4_1 _4646_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ),
    .S0(net387),
    .S1(net376),
    .X(_2286_));
 sky130_fd_sc_hd__mux4_1 _4647_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ),
    .S0(net387),
    .S1(net376),
    .X(_2287_));
 sky130_fd_sc_hd__mux2_1 _4648_ (.A0(_2286_),
    .A1(_2287_),
    .S(net370),
    .X(_2288_));
 sky130_fd_sc_hd__mux4_1 _4649_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ),
    .S0(net387),
    .S1(net376),
    .X(_2289_));
 sky130_fd_sc_hd__mux4_1 _4650_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ),
    .S0(net387),
    .S1(net376),
    .X(_2290_));
 sky130_fd_sc_hd__mux2_1 _4651_ (.A0(_2290_),
    .A1(_2289_),
    .S(net370),
    .X(_2291_));
 sky130_fd_sc_hd__mux2_1 _4652_ (.A0(_2291_),
    .A1(_2288_),
    .S(net368),
    .X(_0009_));
 sky130_fd_sc_hd__mux4_1 _4653_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ),
    .S0(net389),
    .S1(net378),
    .X(_2292_));
 sky130_fd_sc_hd__mux4_1 _4654_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ),
    .S0(net389),
    .S1(net378),
    .X(_2293_));
 sky130_fd_sc_hd__mux2_1 _4655_ (.A0(_2292_),
    .A1(_2293_),
    .S(net370),
    .X(_2294_));
 sky130_fd_sc_hd__mux4_1 _4656_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ),
    .S0(net389),
    .S1(net378),
    .X(_2295_));
 sky130_fd_sc_hd__mux4_1 _4657_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ),
    .S0(net389),
    .S1(net378),
    .X(_2296_));
 sky130_fd_sc_hd__mux2_1 _4658_ (.A0(_2296_),
    .A1(_2295_),
    .S(net370),
    .X(_2297_));
 sky130_fd_sc_hd__mux2_1 _4659_ (.A0(_2297_),
    .A1(_2294_),
    .S(net368),
    .X(_0010_));
 sky130_fd_sc_hd__mux4_1 _4660_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ),
    .S0(net387),
    .S1(net376),
    .X(_2298_));
 sky130_fd_sc_hd__mux4_1 _4661_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ),
    .S0(net387),
    .S1(net376),
    .X(_2299_));
 sky130_fd_sc_hd__mux2_1 _4662_ (.A0(_2298_),
    .A1(_2299_),
    .S(net370),
    .X(_2300_));
 sky130_fd_sc_hd__mux4_1 _4663_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ),
    .S0(net387),
    .S1(net376),
    .X(_2301_));
 sky130_fd_sc_hd__mux4_1 _4664_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ),
    .S0(net387),
    .S1(net376),
    .X(_2302_));
 sky130_fd_sc_hd__mux2_1 _4665_ (.A0(_2302_),
    .A1(_2301_),
    .S(net370),
    .X(_2303_));
 sky130_fd_sc_hd__mux2_1 _4666_ (.A0(_2303_),
    .A1(_2300_),
    .S(net368),
    .X(_0012_));
 sky130_fd_sc_hd__mux4_1 _4667_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ),
    .S0(net392),
    .S1(net381),
    .X(_2304_));
 sky130_fd_sc_hd__mux4_1 _4668_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ),
    .S0(net392),
    .S1(net381),
    .X(_2305_));
 sky130_fd_sc_hd__mux2_1 _4669_ (.A0(_2304_),
    .A1(_2305_),
    .S(net373),
    .X(_2306_));
 sky130_fd_sc_hd__mux4_1 _4670_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ),
    .S0(net392),
    .S1(net381),
    .X(_2307_));
 sky130_fd_sc_hd__mux4_1 _4671_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ),
    .S0(net392),
    .S1(net381),
    .X(_2308_));
 sky130_fd_sc_hd__mux2_1 _4672_ (.A0(_2308_),
    .A1(_2307_),
    .S(net373),
    .X(_2309_));
 sky130_fd_sc_hd__mux2_1 _4673_ (.A0(_2309_),
    .A1(_2306_),
    .S(net369),
    .X(_0013_));
 sky130_fd_sc_hd__mux4_1 _4674_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ),
    .S0(net390),
    .S1(net379),
    .X(_2310_));
 sky130_fd_sc_hd__mux4_1 _4675_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ),
    .S0(net390),
    .S1(net379),
    .X(_2311_));
 sky130_fd_sc_hd__mux2_1 _4676_ (.A0(_2310_),
    .A1(_2311_),
    .S(net371),
    .X(_2312_));
 sky130_fd_sc_hd__mux4_1 _4677_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ),
    .S0(net387),
    .S1(net376),
    .X(_2313_));
 sky130_fd_sc_hd__mux4_1 _4678_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ),
    .S0(net387),
    .S1(net376),
    .X(_2314_));
 sky130_fd_sc_hd__mux2_1 _4679_ (.A0(_2314_),
    .A1(_2313_),
    .S(net371),
    .X(_2315_));
 sky130_fd_sc_hd__mux2_1 _4680_ (.A0(_2315_),
    .A1(_2312_),
    .S(net368),
    .X(_0014_));
 sky130_fd_sc_hd__mux4_1 _4681_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ),
    .S0(net388),
    .S1(net377),
    .X(_2316_));
 sky130_fd_sc_hd__mux4_1 _4682_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ),
    .S0(net388),
    .S1(net377),
    .X(_2317_));
 sky130_fd_sc_hd__mux2_1 _4683_ (.A0(_2316_),
    .A1(_2317_),
    .S(net370),
    .X(_2318_));
 sky130_fd_sc_hd__mux4_1 _4684_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ),
    .S0(net388),
    .S1(net377),
    .X(_2319_));
 sky130_fd_sc_hd__mux4_1 _4685_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ),
    .S0(net388),
    .S1(net377),
    .X(_2320_));
 sky130_fd_sc_hd__mux2_1 _4686_ (.A0(_2320_),
    .A1(_2319_),
    .S(net370),
    .X(_2321_));
 sky130_fd_sc_hd__mux2_1 _4687_ (.A0(_2321_),
    .A1(_2318_),
    .S(net368),
    .X(_0015_));
 sky130_fd_sc_hd__mux4_1 _4688_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ),
    .S0(net391),
    .S1(net380),
    .X(_2322_));
 sky130_fd_sc_hd__mux4_1 _4689_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ),
    .S0(net391),
    .S1(net380),
    .X(_2323_));
 sky130_fd_sc_hd__mux2_1 _4690_ (.A0(_2322_),
    .A1(_2323_),
    .S(net372),
    .X(_2324_));
 sky130_fd_sc_hd__mux4_1 _4691_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ),
    .S0(net391),
    .S1(net380),
    .X(_2325_));
 sky130_fd_sc_hd__mux4_1 _4692_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ),
    .S0(net391),
    .S1(net380),
    .X(_2326_));
 sky130_fd_sc_hd__mux2_1 _4693_ (.A0(_2326_),
    .A1(_2325_),
    .S(net372),
    .X(_2327_));
 sky130_fd_sc_hd__mux2_1 _4694_ (.A0(_2327_),
    .A1(_2324_),
    .S(net368),
    .X(_0016_));
 sky130_fd_sc_hd__mux4_1 _4695_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ),
    .S0(net393),
    .S1(net381),
    .X(_2328_));
 sky130_fd_sc_hd__mux4_1 _4696_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ),
    .S0(net392),
    .S1(net381),
    .X(_2329_));
 sky130_fd_sc_hd__mux2_1 _4697_ (.A0(_2328_),
    .A1(_2329_),
    .S(net373),
    .X(_2330_));
 sky130_fd_sc_hd__mux4_1 _4698_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ),
    .S0(net389),
    .S1(net378),
    .X(_2331_));
 sky130_fd_sc_hd__mux4_1 _4699_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ),
    .S0(net389),
    .S1(net378),
    .X(_2332_));
 sky130_fd_sc_hd__mux2_1 _4700_ (.A0(_2332_),
    .A1(_2331_),
    .S(net371),
    .X(_2333_));
 sky130_fd_sc_hd__mux2_1 _4701_ (.A0(_2333_),
    .A1(_2330_),
    .S(net368),
    .X(_0017_));
 sky130_fd_sc_hd__mux4_1 _4702_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ),
    .S0(net388),
    .S1(net377),
    .X(_2334_));
 sky130_fd_sc_hd__mux4_1 _4703_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ),
    .S0(net388),
    .S1(net376),
    .X(_2335_));
 sky130_fd_sc_hd__mux2_1 _4704_ (.A0(_2334_),
    .A1(_2335_),
    .S(net370),
    .X(_2336_));
 sky130_fd_sc_hd__mux4_1 _4705_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ),
    .S0(net387),
    .S1(net377),
    .X(_2337_));
 sky130_fd_sc_hd__mux4_1 _4706_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ),
    .S0(net387),
    .S1(net377),
    .X(_2338_));
 sky130_fd_sc_hd__mux2_1 _4707_ (.A0(_2338_),
    .A1(_2337_),
    .S(net370),
    .X(_2339_));
 sky130_fd_sc_hd__mux2_1 _4708_ (.A0(_2339_),
    .A1(_2336_),
    .S(net368),
    .X(_0018_));
 sky130_fd_sc_hd__mux4_1 _4709_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ),
    .S0(net388),
    .S1(net377),
    .X(_2340_));
 sky130_fd_sc_hd__mux4_1 _4710_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ),
    .S0(net388),
    .S1(net377),
    .X(_2341_));
 sky130_fd_sc_hd__mux2_1 _4711_ (.A0(_2340_),
    .A1(_2341_),
    .S(net370),
    .X(_2342_));
 sky130_fd_sc_hd__mux4_1 _4712_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ),
    .S0(net391),
    .S1(net380),
    .X(_2343_));
 sky130_fd_sc_hd__mux4_1 _4713_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ),
    .S0(net391),
    .S1(net380),
    .X(_2344_));
 sky130_fd_sc_hd__mux2_1 _4714_ (.A0(_2344_),
    .A1(_2343_),
    .S(net372),
    .X(_2345_));
 sky130_fd_sc_hd__mux2_1 _4715_ (.A0(_2345_),
    .A1(_2342_),
    .S(net368),
    .X(_0019_));
 sky130_fd_sc_hd__mux4_1 _4716_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ),
    .S0(net390),
    .S1(net379),
    .X(_2346_));
 sky130_fd_sc_hd__mux4_1 _4717_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ),
    .S0(net390),
    .S1(net378),
    .X(_2347_));
 sky130_fd_sc_hd__mux2_1 _4718_ (.A0(_2346_),
    .A1(_2347_),
    .S(net371),
    .X(_2348_));
 sky130_fd_sc_hd__mux4_1 _4719_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ),
    .S0(net390),
    .S1(net379),
    .X(_2349_));
 sky130_fd_sc_hd__mux4_1 _4720_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ),
    .S0(net390),
    .S1(net379),
    .X(_2350_));
 sky130_fd_sc_hd__mux2_1 _4721_ (.A0(_2350_),
    .A1(_2349_),
    .S(net371),
    .X(_2351_));
 sky130_fd_sc_hd__mux2_1 _4722_ (.A0(_2351_),
    .A1(_2348_),
    .S(net368),
    .X(_0020_));
 sky130_fd_sc_hd__mux4_1 _4723_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ),
    .S0(net391),
    .S1(net380),
    .X(_2352_));
 sky130_fd_sc_hd__mux4_1 _4724_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ),
    .S0(net391),
    .S1(net380),
    .X(_2353_));
 sky130_fd_sc_hd__mux2_1 _4725_ (.A0(_2352_),
    .A1(_2353_),
    .S(net372),
    .X(_2354_));
 sky130_fd_sc_hd__mux4_1 _4726_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ),
    .S0(net391),
    .S1(net380),
    .X(_2355_));
 sky130_fd_sc_hd__mux4_1 _4727_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ),
    .S0(net391),
    .S1(net380),
    .X(_2356_));
 sky130_fd_sc_hd__mux2_1 _4728_ (.A0(_2356_),
    .A1(_2355_),
    .S(net372),
    .X(_2357_));
 sky130_fd_sc_hd__mux2_1 _4729_ (.A0(_2357_),
    .A1(_2354_),
    .S(net368),
    .X(_0021_));
 sky130_fd_sc_hd__mux4_1 _4730_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ),
    .S0(net389),
    .S1(net378),
    .X(_2358_));
 sky130_fd_sc_hd__mux4_1 _4731_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ),
    .S0(net389),
    .S1(net378),
    .X(_2359_));
 sky130_fd_sc_hd__mux2_1 _4732_ (.A0(_2358_),
    .A1(_2359_),
    .S(net370),
    .X(_2360_));
 sky130_fd_sc_hd__mux4_1 _4733_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ),
    .S0(net388),
    .S1(net376),
    .X(_2361_));
 sky130_fd_sc_hd__mux4_1 _4734_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ),
    .S0(net388),
    .S1(net377),
    .X(_2362_));
 sky130_fd_sc_hd__mux2_1 _4735_ (.A0(_2362_),
    .A1(_2361_),
    .S(net371),
    .X(_2363_));
 sky130_fd_sc_hd__mux2_1 _4736_ (.A0(_2363_),
    .A1(_2360_),
    .S(net368),
    .X(_0023_));
 sky130_fd_sc_hd__mux4_1 _4737_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ),
    .S0(net393),
    .S1(net384),
    .X(_2364_));
 sky130_fd_sc_hd__mux4_1 _4738_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ),
    .S0(net393),
    .S1(net386),
    .X(_2365_));
 sky130_fd_sc_hd__mux2_1 _4739_ (.A0(_2364_),
    .A1(_2365_),
    .S(net373),
    .X(_2366_));
 sky130_fd_sc_hd__mux4_1 _4740_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ),
    .S0(net393),
    .S1(net381),
    .X(_2367_));
 sky130_fd_sc_hd__mux4_1 _4741_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ),
    .S0(net393),
    .S1(net379),
    .X(_2368_));
 sky130_fd_sc_hd__mux2_1 _4742_ (.A0(_2368_),
    .A1(_2367_),
    .S(net373),
    .X(_2369_));
 sky130_fd_sc_hd__mux2_1 _4743_ (.A0(_2369_),
    .A1(_2366_),
    .S(net369),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _4744_ (.A(net453),
    .B(net1410),
    .X(_0069_));
 sky130_fd_sc_hd__and2_1 _4745_ (.A(net453),
    .B(net1996),
    .X(_0080_));
 sky130_fd_sc_hd__and2_1 _4746_ (.A(net446),
    .B(net923),
    .X(_0091_));
 sky130_fd_sc_hd__and2_1 _4747_ (.A(net446),
    .B(net610),
    .X(_0094_));
 sky130_fd_sc_hd__and2_1 _4748_ (.A(net439),
    .B(net2173),
    .X(_0095_));
 sky130_fd_sc_hd__and2_1 _4749_ (.A(net445),
    .B(net660),
    .X(_0096_));
 sky130_fd_sc_hd__and2_1 _4750_ (.A(net448),
    .B(net1558),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _4751_ (.A(net452),
    .B(net1017),
    .X(_0098_));
 sky130_fd_sc_hd__and2_1 _4752_ (.A(net451),
    .B(net2133),
    .X(_0099_));
 sky130_fd_sc_hd__and2_1 _4753_ (.A(net453),
    .B(net2191),
    .X(_0100_));
 sky130_fd_sc_hd__and2_1 _4754_ (.A(net453),
    .B(net2033),
    .X(_0070_));
 sky130_fd_sc_hd__and2_1 _4755_ (.A(net434),
    .B(net2071),
    .X(_0071_));
 sky130_fd_sc_hd__and2_1 _4756_ (.A(net453),
    .B(net2137),
    .X(_0072_));
 sky130_fd_sc_hd__and2_1 _4757_ (.A(net453),
    .B(net1970),
    .X(_0073_));
 sky130_fd_sc_hd__and2_1 _4758_ (.A(net446),
    .B(net2066),
    .X(_0074_));
 sky130_fd_sc_hd__and2_1 _4759_ (.A(net433),
    .B(net2174),
    .X(_0075_));
 sky130_fd_sc_hd__and2_1 _4760_ (.A(net434),
    .B(net2104),
    .X(_0076_));
 sky130_fd_sc_hd__and2_1 _4761_ (.A(net455),
    .B(net2007),
    .X(_0077_));
 sky130_fd_sc_hd__and2_1 _4762_ (.A(net443),
    .B(net1897),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _4763_ (.A(net432),
    .B(net2113),
    .X(_0079_));
 sky130_fd_sc_hd__and2_1 _4764_ (.A(net429),
    .B(net2045),
    .X(_0081_));
 sky130_fd_sc_hd__and2_1 _4765_ (.A(net444),
    .B(net2099),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _4766_ (.A(net443),
    .B(net2037),
    .X(_0083_));
 sky130_fd_sc_hd__and2_1 _4767_ (.A(net436),
    .B(net2092),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _4768_ (.A(net439),
    .B(net2016),
    .X(_0085_));
 sky130_fd_sc_hd__and2_1 _4769_ (.A(net434),
    .B(net2105),
    .X(_0086_));
 sky130_fd_sc_hd__and2_1 _4770_ (.A(net440),
    .B(net2190),
    .X(_0087_));
 sky130_fd_sc_hd__and2_1 _4771_ (.A(net439),
    .B(net2035),
    .X(_0088_));
 sky130_fd_sc_hd__and2_1 _4772_ (.A(net441),
    .B(net2253),
    .X(_0089_));
 sky130_fd_sc_hd__and2_1 _4773_ (.A(net442),
    .B(net2077),
    .X(_0090_));
 sky130_fd_sc_hd__and2_1 _4774_ (.A(net434),
    .B(net2076),
    .X(_0092_));
 sky130_fd_sc_hd__and2_1 _4775_ (.A(net459),
    .B(net2167),
    .X(_0093_));
 sky130_fd_sc_hd__mux4_1 _4776_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ),
    .S0(net424),
    .S1(net414),
    .X(_2370_));
 sky130_fd_sc_hd__mux4_1 _4777_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ),
    .S0(net424),
    .S1(net414),
    .X(_2371_));
 sky130_fd_sc_hd__mux2_1 _4778_ (.A0(_2370_),
    .A1(_2371_),
    .S(net404),
    .X(_2372_));
 sky130_fd_sc_hd__mux4_1 _4779_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ),
    .S0(net424),
    .S1(net414),
    .X(_2373_));
 sky130_fd_sc_hd__mux4_1 _4780_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ),
    .S0(net424),
    .S1(net414),
    .X(_2374_));
 sky130_fd_sc_hd__mux2_1 _4781_ (.A0(_2374_),
    .A1(_2373_),
    .S(net404),
    .X(_2375_));
 sky130_fd_sc_hd__mux2_1 _4782_ (.A0(_2375_),
    .A1(_2372_),
    .S(net398),
    .X(_0032_));
 sky130_fd_sc_hd__mux4_1 _4783_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ),
    .S0(net424),
    .S1(net414),
    .X(_2376_));
 sky130_fd_sc_hd__mux4_1 _4784_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ),
    .S0(net424),
    .S1(net414),
    .X(_2377_));
 sky130_fd_sc_hd__mux2_1 _4785_ (.A0(_2376_),
    .A1(_2377_),
    .S(net404),
    .X(_2378_));
 sky130_fd_sc_hd__mux4_1 _4786_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ),
    .S0(net424),
    .S1(net414),
    .X(_2379_));
 sky130_fd_sc_hd__mux4_1 _4787_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ),
    .S0(net424),
    .S1(net414),
    .X(_2380_));
 sky130_fd_sc_hd__mux2_1 _4788_ (.A0(_2380_),
    .A1(_2379_),
    .S(net404),
    .X(_2381_));
 sky130_fd_sc_hd__mux2_1 _4789_ (.A0(_2381_),
    .A1(_2378_),
    .S(net398),
    .X(_0043_));
 sky130_fd_sc_hd__mux4_1 _4790_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ),
    .S0(net422),
    .S1(net413),
    .X(_2382_));
 sky130_fd_sc_hd__mux4_1 _4791_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ),
    .S0(net422),
    .S1(net413),
    .X(_2383_));
 sky130_fd_sc_hd__mux2_1 _4792_ (.A0(_2382_),
    .A1(_2383_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ),
    .X(_2384_));
 sky130_fd_sc_hd__mux4_1 _4793_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ),
    .S0(net424),
    .S1(net412),
    .X(_2385_));
 sky130_fd_sc_hd__mux4_1 _4794_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ),
    .S0(net424),
    .S1(net413),
    .X(_2386_));
 sky130_fd_sc_hd__mux2_1 _4795_ (.A0(_2386_),
    .A1(_2385_),
    .S(net404),
    .X(_2387_));
 sky130_fd_sc_hd__mux2_1 _4796_ (.A0(_2387_),
    .A1(_2384_),
    .S(net398),
    .X(_0054_));
 sky130_fd_sc_hd__mux4_1 _4797_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ),
    .S0(net423),
    .S1(net413),
    .X(_2388_));
 sky130_fd_sc_hd__mux4_1 _4798_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ),
    .S0(net423),
    .S1(net412),
    .X(_2389_));
 sky130_fd_sc_hd__mux2_1 _4799_ (.A0(_2388_),
    .A1(_2389_),
    .S(net403),
    .X(_2390_));
 sky130_fd_sc_hd__mux4_1 _4800_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ),
    .S0(net422),
    .S1(net413),
    .X(_2391_));
 sky130_fd_sc_hd__mux4_1 _4801_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ),
    .S0(net423),
    .S1(net413),
    .X(_2392_));
 sky130_fd_sc_hd__mux2_1 _4802_ (.A0(_2392_),
    .A1(_2391_),
    .S(net403),
    .X(_2393_));
 sky130_fd_sc_hd__mux2_1 _4803_ (.A0(_2393_),
    .A1(_2390_),
    .S(net398),
    .X(_0057_));
 sky130_fd_sc_hd__mux4_1 _4804_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ),
    .S0(net418),
    .S1(net409),
    .X(_2394_));
 sky130_fd_sc_hd__mux4_1 _4805_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ),
    .S0(net418),
    .S1(net409),
    .X(_2395_));
 sky130_fd_sc_hd__mux2_1 _4806_ (.A0(_2394_),
    .A1(_2395_),
    .S(net402),
    .X(_2396_));
 sky130_fd_sc_hd__mux4_1 _4807_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ),
    .S0(net418),
    .S1(net409),
    .X(_2397_));
 sky130_fd_sc_hd__mux4_1 _4808_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ),
    .S0(net418),
    .S1(net409),
    .X(_2398_));
 sky130_fd_sc_hd__mux2_1 _4809_ (.A0(_2398_),
    .A1(_2397_),
    .S(net402),
    .X(_2399_));
 sky130_fd_sc_hd__mux2_1 _4810_ (.A0(_2399_),
    .A1(_2396_),
    .S(net397),
    .X(_0058_));
 sky130_fd_sc_hd__mux4_1 _4811_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ),
    .S0(net420),
    .S1(net410),
    .X(_2400_));
 sky130_fd_sc_hd__mux4_1 _4812_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ),
    .S0(net420),
    .S1(net410),
    .X(_2401_));
 sky130_fd_sc_hd__mux2_1 _4813_ (.A0(_2400_),
    .A1(_2401_),
    .S(net403),
    .X(_2402_));
 sky130_fd_sc_hd__mux4_1 _4814_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ),
    .S0(net420),
    .S1(net410),
    .X(_2403_));
 sky130_fd_sc_hd__mux4_1 _4815_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ),
    .S0(net420),
    .S1(net410),
    .X(_2404_));
 sky130_fd_sc_hd__mux2_1 _4816_ (.A0(_2404_),
    .A1(_2403_),
    .S(net403),
    .X(_2405_));
 sky130_fd_sc_hd__mux2_1 _4817_ (.A0(_2405_),
    .A1(_2402_),
    .S(net398),
    .X(_0059_));
 sky130_fd_sc_hd__mux4_1 _4818_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ),
    .S0(net422),
    .S1(net412),
    .X(_2406_));
 sky130_fd_sc_hd__mux4_1 _4819_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ),
    .S0(net422),
    .S1(net412),
    .X(_2407_));
 sky130_fd_sc_hd__mux2_1 _4820_ (.A0(_2406_),
    .A1(_2407_),
    .S(net404),
    .X(_2408_));
 sky130_fd_sc_hd__mux4_1 _4821_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ),
    .S0(net422),
    .S1(net412),
    .X(_2409_));
 sky130_fd_sc_hd__mux4_1 _4822_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ),
    .S0(net422),
    .S1(net412),
    .X(_2410_));
 sky130_fd_sc_hd__mux2_1 _4823_ (.A0(_2410_),
    .A1(_2409_),
    .S(net404),
    .X(_2411_));
 sky130_fd_sc_hd__mux2_1 _4824_ (.A0(_2411_),
    .A1(_2408_),
    .S(net398),
    .X(_0060_));
 sky130_fd_sc_hd__mux4_1 _4825_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ),
    .S0(net418),
    .S1(net408),
    .X(_2412_));
 sky130_fd_sc_hd__mux4_1 _4826_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ),
    .S0(net419),
    .S1(net408),
    .X(_2413_));
 sky130_fd_sc_hd__mux2_1 _4827_ (.A0(_2412_),
    .A1(_2413_),
    .S(net402),
    .X(_2414_));
 sky130_fd_sc_hd__mux4_1 _4828_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ),
    .S0(net419),
    .S1(net409),
    .X(_2415_));
 sky130_fd_sc_hd__mux4_1 _4829_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ),
    .S0(net419),
    .S1(net409),
    .X(_2416_));
 sky130_fd_sc_hd__mux2_1 _4830_ (.A0(_2416_),
    .A1(_2415_),
    .S(net402),
    .X(_2417_));
 sky130_fd_sc_hd__mux2_1 _4831_ (.A0(_2417_),
    .A1(_2414_),
    .S(net397),
    .X(_0061_));
 sky130_fd_sc_hd__mux4_1 _4832_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ),
    .S0(net424),
    .S1(net414),
    .X(_2418_));
 sky130_fd_sc_hd__mux4_1 _4833_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ),
    .S0(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .S1(net414),
    .X(_2419_));
 sky130_fd_sc_hd__mux2_1 _4834_ (.A0(_2418_),
    .A1(_2419_),
    .S(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ),
    .X(_2420_));
 sky130_fd_sc_hd__mux4_1 _4835_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ),
    .S0(net424),
    .S1(net414),
    .X(_2421_));
 sky130_fd_sc_hd__mux4_1 _4836_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ),
    .S0(net424),
    .S1(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ),
    .X(_2422_));
 sky130_fd_sc_hd__mux2_1 _4837_ (.A0(_2422_),
    .A1(_2421_),
    .S(net404),
    .X(_2423_));
 sky130_fd_sc_hd__mux2_1 _4838_ (.A0(_2423_),
    .A1(_2420_),
    .S(net398),
    .X(_0062_));
 sky130_fd_sc_hd__mux4_1 _4839_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ),
    .S0(net422),
    .S1(net412),
    .X(_2424_));
 sky130_fd_sc_hd__mux4_1 _4840_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ),
    .S0(net422),
    .S1(net412),
    .X(_2425_));
 sky130_fd_sc_hd__mux2_1 _4841_ (.A0(_2424_),
    .A1(_2425_),
    .S(net404),
    .X(_2426_));
 sky130_fd_sc_hd__mux4_1 _4842_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ),
    .S0(net422),
    .S1(net412),
    .X(_2427_));
 sky130_fd_sc_hd__mux4_1 _4843_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ),
    .S0(net422),
    .S1(net412),
    .X(_2428_));
 sky130_fd_sc_hd__mux2_1 _4844_ (.A0(_2428_),
    .A1(_2427_),
    .S(net403),
    .X(_2429_));
 sky130_fd_sc_hd__mux2_1 _4845_ (.A0(_2429_),
    .A1(_2426_),
    .S(net398),
    .X(_0063_));
 sky130_fd_sc_hd__mux4_1 _4846_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ),
    .S0(net422),
    .S1(net412),
    .X(_2430_));
 sky130_fd_sc_hd__mux4_1 _4847_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ),
    .S0(net422),
    .S1(net412),
    .X(_2431_));
 sky130_fd_sc_hd__mux2_1 _4848_ (.A0(_2430_),
    .A1(_2431_),
    .S(net404),
    .X(_2432_));
 sky130_fd_sc_hd__mux4_1 _4849_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ),
    .S0(net422),
    .S1(net412),
    .X(_2433_));
 sky130_fd_sc_hd__mux4_1 _4850_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ),
    .S0(net422),
    .S1(net412),
    .X(_2434_));
 sky130_fd_sc_hd__mux2_1 _4851_ (.A0(_2434_),
    .A1(_2433_),
    .S(net404),
    .X(_2435_));
 sky130_fd_sc_hd__mux2_1 _4852_ (.A0(_2435_),
    .A1(_2432_),
    .S(net398),
    .X(_0033_));
 sky130_fd_sc_hd__mux4_1 _4853_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ),
    .S0(net417),
    .S1(net407),
    .X(_2436_));
 sky130_fd_sc_hd__mux4_1 _4854_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ),
    .S0(net417),
    .S1(net407),
    .X(_2437_));
 sky130_fd_sc_hd__mux2_1 _4855_ (.A0(_2436_),
    .A1(_2437_),
    .S(net401),
    .X(_2438_));
 sky130_fd_sc_hd__mux4_1 _4856_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ),
    .S0(net417),
    .S1(net407),
    .X(_2439_));
 sky130_fd_sc_hd__mux4_1 _4857_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ),
    .S0(net417),
    .S1(net407),
    .X(_2440_));
 sky130_fd_sc_hd__mux2_1 _4858_ (.A0(_2440_),
    .A1(_2439_),
    .S(net401),
    .X(_2441_));
 sky130_fd_sc_hd__mux2_1 _4859_ (.A0(_2441_),
    .A1(_2438_),
    .S(net397),
    .X(_0034_));
 sky130_fd_sc_hd__mux4_1 _4860_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ),
    .S0(net423),
    .S1(net413),
    .X(_2442_));
 sky130_fd_sc_hd__mux4_1 _4861_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ),
    .S0(net423),
    .S1(net413),
    .X(_2443_));
 sky130_fd_sc_hd__mux2_1 _4862_ (.A0(_2442_),
    .A1(_2443_),
    .S(net404),
    .X(_2444_));
 sky130_fd_sc_hd__mux4_1 _4863_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ),
    .S0(net423),
    .S1(net413),
    .X(_2445_));
 sky130_fd_sc_hd__mux4_1 _4864_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ),
    .S0(net423),
    .S1(net413),
    .X(_2446_));
 sky130_fd_sc_hd__mux2_1 _4865_ (.A0(_2446_),
    .A1(_2445_),
    .S(net403),
    .X(_2447_));
 sky130_fd_sc_hd__mux2_1 _4866_ (.A0(_2447_),
    .A1(_2444_),
    .S(net398),
    .X(_0035_));
 sky130_fd_sc_hd__mux4_1 _4867_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ),
    .S0(net423),
    .S1(net413),
    .X(_2448_));
 sky130_fd_sc_hd__mux4_1 _4868_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ),
    .S0(net421),
    .S1(net411),
    .X(_2449_));
 sky130_fd_sc_hd__mux2_1 _4869_ (.A0(_2448_),
    .A1(_2449_),
    .S(net403),
    .X(_2450_));
 sky130_fd_sc_hd__mux4_1 _4870_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ),
    .S0(net421),
    .S1(net411),
    .X(_2451_));
 sky130_fd_sc_hd__mux4_1 _4871_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ),
    .S0(net421),
    .S1(net411),
    .X(_2452_));
 sky130_fd_sc_hd__mux2_1 _4872_ (.A0(_2452_),
    .A1(_2451_),
    .S(net403),
    .X(_2453_));
 sky130_fd_sc_hd__mux2_1 _4873_ (.A0(_2453_),
    .A1(_2450_),
    .S(net398),
    .X(_0036_));
 sky130_fd_sc_hd__mux4_1 _4874_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ),
    .S0(net420),
    .S1(net410),
    .X(_2454_));
 sky130_fd_sc_hd__mux4_1 _4875_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ),
    .S0(net421),
    .S1(net410),
    .X(_2455_));
 sky130_fd_sc_hd__mux2_1 _4876_ (.A0(_2454_),
    .A1(_2455_),
    .S(net403),
    .X(_2456_));
 sky130_fd_sc_hd__mux4_1 _4877_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ),
    .S0(net420),
    .S1(net410),
    .X(_2457_));
 sky130_fd_sc_hd__mux4_1 _4878_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ),
    .S0(net420),
    .S1(net410),
    .X(_2458_));
 sky130_fd_sc_hd__mux2_1 _4879_ (.A0(_2458_),
    .A1(_2457_),
    .S(net403),
    .X(_2459_));
 sky130_fd_sc_hd__mux2_1 _4880_ (.A0(_2459_),
    .A1(_2456_),
    .S(net398),
    .X(_0037_));
 sky130_fd_sc_hd__mux4_1 _4881_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ),
    .S0(net415),
    .S1(net405),
    .X(_2460_));
 sky130_fd_sc_hd__mux4_1 _4882_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ),
    .S0(net415),
    .S1(net405),
    .X(_2461_));
 sky130_fd_sc_hd__mux2_1 _4883_ (.A0(_2460_),
    .A1(_2461_),
    .S(net400),
    .X(_2462_));
 sky130_fd_sc_hd__mux4_1 _4884_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ),
    .S0(net415),
    .S1(net405),
    .X(_2463_));
 sky130_fd_sc_hd__mux4_1 _4885_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ),
    .S0(net415),
    .S1(net405),
    .X(_2464_));
 sky130_fd_sc_hd__mux2_1 _4886_ (.A0(_2464_),
    .A1(_2463_),
    .S(net400),
    .X(_2465_));
 sky130_fd_sc_hd__mux2_1 _4887_ (.A0(_2465_),
    .A1(_2462_),
    .S(net397),
    .X(_0038_));
 sky130_fd_sc_hd__mux4_1 _4888_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ),
    .S0(net417),
    .S1(net407),
    .X(_2466_));
 sky130_fd_sc_hd__mux4_1 _4889_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ),
    .S0(net420),
    .S1(net410),
    .X(_2467_));
 sky130_fd_sc_hd__mux2_1 _4890_ (.A0(_2466_),
    .A1(_2467_),
    .S(net400),
    .X(_2468_));
 sky130_fd_sc_hd__mux4_1 _4891_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ),
    .S0(net420),
    .S1(net410),
    .X(_2469_));
 sky130_fd_sc_hd__mux4_1 _4892_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ),
    .S0(net417),
    .S1(net407),
    .X(_2470_));
 sky130_fd_sc_hd__mux2_1 _4893_ (.A0(_2470_),
    .A1(_2469_),
    .S(net400),
    .X(_2471_));
 sky130_fd_sc_hd__mux2_1 _4894_ (.A0(_2471_),
    .A1(_2468_),
    .S(net397),
    .X(_0039_));
 sky130_fd_sc_hd__mux4_1 _4895_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ),
    .S0(net422),
    .S1(net412),
    .X(_2472_));
 sky130_fd_sc_hd__mux4_1 _4896_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ),
    .S0(net423),
    .S1(net412),
    .X(_2473_));
 sky130_fd_sc_hd__mux2_1 _4897_ (.A0(_2472_),
    .A1(_2473_),
    .S(net403),
    .X(_2474_));
 sky130_fd_sc_hd__mux4_1 _4898_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ),
    .S0(net420),
    .S1(net411),
    .X(_2475_));
 sky130_fd_sc_hd__mux4_1 _4899_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ),
    .S0(net421),
    .S1(net410),
    .X(_2476_));
 sky130_fd_sc_hd__mux2_1 _4900_ (.A0(_2476_),
    .A1(_2475_),
    .S(net403),
    .X(_2477_));
 sky130_fd_sc_hd__mux2_1 _4901_ (.A0(_2477_),
    .A1(_2474_),
    .S(net398),
    .X(_0040_));
 sky130_fd_sc_hd__mux4_1 _4902_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ),
    .S0(net415),
    .S1(net405),
    .X(_2478_));
 sky130_fd_sc_hd__mux4_1 _4903_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ),
    .S0(net415),
    .S1(net405),
    .X(_2479_));
 sky130_fd_sc_hd__mux2_1 _4904_ (.A0(_2478_),
    .A1(_2479_),
    .S(net400),
    .X(_2480_));
 sky130_fd_sc_hd__mux4_1 _4905_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ),
    .S0(net415),
    .S1(net405),
    .X(_2481_));
 sky130_fd_sc_hd__mux4_1 _4906_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ),
    .S0(net415),
    .S1(net405),
    .X(_2482_));
 sky130_fd_sc_hd__mux2_1 _4907_ (.A0(_2482_),
    .A1(_2481_),
    .S(net400),
    .X(_2483_));
 sky130_fd_sc_hd__mux2_1 _4908_ (.A0(_2483_),
    .A1(_2480_),
    .S(net397),
    .X(_0041_));
 sky130_fd_sc_hd__mux4_1 _4909_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ),
    .S0(net417),
    .S1(net407),
    .X(_2484_));
 sky130_fd_sc_hd__mux4_1 _4910_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ),
    .S0(net417),
    .S1(net407),
    .X(_2485_));
 sky130_fd_sc_hd__mux2_1 _4911_ (.A0(_2484_),
    .A1(_2485_),
    .S(net401),
    .X(_2486_));
 sky130_fd_sc_hd__mux4_1 _4912_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ),
    .S0(net417),
    .S1(net407),
    .X(_2487_));
 sky130_fd_sc_hd__mux4_1 _4913_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ),
    .S0(net417),
    .S1(net407),
    .X(_2488_));
 sky130_fd_sc_hd__mux2_1 _4914_ (.A0(_2488_),
    .A1(_2487_),
    .S(net400),
    .X(_2489_));
 sky130_fd_sc_hd__mux2_1 _4915_ (.A0(_2489_),
    .A1(_2486_),
    .S(net397),
    .X(_0042_));
 sky130_fd_sc_hd__mux4_1 _4916_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ),
    .S0(net415),
    .S1(net405),
    .X(_2490_));
 sky130_fd_sc_hd__mux4_1 _4917_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ),
    .S0(net415),
    .S1(net405),
    .X(_2491_));
 sky130_fd_sc_hd__mux2_1 _4918_ (.A0(_2490_),
    .A1(_2491_),
    .S(net400),
    .X(_2492_));
 sky130_fd_sc_hd__mux4_1 _4919_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ),
    .S0(net415),
    .S1(net405),
    .X(_2493_));
 sky130_fd_sc_hd__mux4_1 _4920_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ),
    .S0(net415),
    .S1(net405),
    .X(_2494_));
 sky130_fd_sc_hd__mux2_1 _4921_ (.A0(_2494_),
    .A1(_2493_),
    .S(net400),
    .X(_2495_));
 sky130_fd_sc_hd__mux2_1 _4922_ (.A0(_2495_),
    .A1(_2492_),
    .S(net397),
    .X(_0044_));
 sky130_fd_sc_hd__mux4_1 _4923_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ),
    .S0(net420),
    .S1(net410),
    .X(_2496_));
 sky130_fd_sc_hd__mux4_1 _4924_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ),
    .S0(net420),
    .S1(net410),
    .X(_2497_));
 sky130_fd_sc_hd__mux2_1 _4925_ (.A0(_2496_),
    .A1(_2497_),
    .S(net403),
    .X(_2498_));
 sky130_fd_sc_hd__mux4_1 _4926_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ),
    .S0(net420),
    .S1(net411),
    .X(_2499_));
 sky130_fd_sc_hd__mux4_1 _4927_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ),
    .S0(net420),
    .S1(net410),
    .X(_2500_));
 sky130_fd_sc_hd__mux2_1 _4928_ (.A0(_2500_),
    .A1(_2499_),
    .S(net403),
    .X(_2501_));
 sky130_fd_sc_hd__mux2_1 _4929_ (.A0(_2501_),
    .A1(_2498_),
    .S(net398),
    .X(_0045_));
 sky130_fd_sc_hd__mux4_1 _4930_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ),
    .S0(net417),
    .S1(net408),
    .X(_2502_));
 sky130_fd_sc_hd__mux4_1 _4931_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ),
    .S0(net417),
    .S1(net407),
    .X(_2503_));
 sky130_fd_sc_hd__mux2_1 _4932_ (.A0(_2502_),
    .A1(_2503_),
    .S(net400),
    .X(_2504_));
 sky130_fd_sc_hd__mux4_1 _4933_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ),
    .S0(net415),
    .S1(net406),
    .X(_2505_));
 sky130_fd_sc_hd__mux4_1 _4934_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ),
    .S0(net418),
    .S1(net406),
    .X(_2506_));
 sky130_fd_sc_hd__mux2_1 _4935_ (.A0(_2506_),
    .A1(_2505_),
    .S(net400),
    .X(_2507_));
 sky130_fd_sc_hd__mux2_1 _4936_ (.A0(_2507_),
    .A1(_2504_),
    .S(net397),
    .X(_0046_));
 sky130_fd_sc_hd__mux4_1 _4937_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ),
    .S0(net416),
    .S1(net406),
    .X(_2508_));
 sky130_fd_sc_hd__mux4_1 _4938_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ),
    .S0(net416),
    .S1(net406),
    .X(_2509_));
 sky130_fd_sc_hd__mux2_1 _4939_ (.A0(_2508_),
    .A1(_2509_),
    .S(net400),
    .X(_2510_));
 sky130_fd_sc_hd__mux4_1 _4940_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ),
    .S0(net416),
    .S1(net405),
    .X(_2511_));
 sky130_fd_sc_hd__mux4_1 _4941_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ),
    .S0(net415),
    .S1(net405),
    .X(_2512_));
 sky130_fd_sc_hd__mux2_1 _4942_ (.A0(_2512_),
    .A1(_2511_),
    .S(net400),
    .X(_2513_));
 sky130_fd_sc_hd__mux2_1 _4943_ (.A0(_2513_),
    .A1(_2510_),
    .S(net397),
    .X(_0047_));
 sky130_fd_sc_hd__mux4_1 _4944_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ),
    .S0(net418),
    .S1(net406),
    .X(_2514_));
 sky130_fd_sc_hd__mux4_1 _4945_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ),
    .S0(net418),
    .S1(net406),
    .X(_2515_));
 sky130_fd_sc_hd__mux2_1 _4946_ (.A0(_2514_),
    .A1(_2515_),
    .S(net402),
    .X(_2516_));
 sky130_fd_sc_hd__mux4_1 _4947_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ),
    .S0(net418),
    .S1(net409),
    .X(_2517_));
 sky130_fd_sc_hd__mux4_1 _4948_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ),
    .S0(net418),
    .S1(net409),
    .X(_2518_));
 sky130_fd_sc_hd__mux2_1 _4949_ (.A0(_2518_),
    .A1(_2517_),
    .S(net402),
    .X(_2519_));
 sky130_fd_sc_hd__mux2_1 _4950_ (.A0(_2519_),
    .A1(_2516_),
    .S(net399),
    .X(_0048_));
 sky130_fd_sc_hd__mux4_1 _4951_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ),
    .S0(net421),
    .S1(net410),
    .X(_2520_));
 sky130_fd_sc_hd__mux4_1 _4952_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ),
    .S0(net420),
    .S1(net410),
    .X(_2521_));
 sky130_fd_sc_hd__mux2_1 _4953_ (.A0(_2520_),
    .A1(_2521_),
    .S(net401),
    .X(_2522_));
 sky130_fd_sc_hd__mux4_1 _4954_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ),
    .S0(net417),
    .S1(net407),
    .X(_2523_));
 sky130_fd_sc_hd__mux4_1 _4955_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ),
    .S0(net417),
    .S1(net407),
    .X(_2524_));
 sky130_fd_sc_hd__mux2_1 _4956_ (.A0(_2524_),
    .A1(_2523_),
    .S(net401),
    .X(_2525_));
 sky130_fd_sc_hd__mux2_1 _4957_ (.A0(_2525_),
    .A1(_2522_),
    .S(net397),
    .X(_0049_));
 sky130_fd_sc_hd__mux4_1 _4958_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ),
    .S0(net415),
    .S1(net406),
    .X(_2526_));
 sky130_fd_sc_hd__mux4_1 _4959_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ),
    .S0(net416),
    .S1(net406),
    .X(_2527_));
 sky130_fd_sc_hd__mux2_1 _4960_ (.A0(_2526_),
    .A1(_2527_),
    .S(net400),
    .X(_2528_));
 sky130_fd_sc_hd__mux4_1 _4961_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ),
    .S0(net416),
    .S1(net406),
    .X(_2529_));
 sky130_fd_sc_hd__mux4_1 _4962_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ),
    .S0(net416),
    .S1(net406),
    .X(_2530_));
 sky130_fd_sc_hd__mux2_1 _4963_ (.A0(_2530_),
    .A1(_2529_),
    .S(net400),
    .X(_2531_));
 sky130_fd_sc_hd__mux2_1 _4964_ (.A0(_2531_),
    .A1(_2528_),
    .S(net397),
    .X(_0050_));
 sky130_fd_sc_hd__mux4_1 _4965_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ),
    .S0(net416),
    .S1(net406),
    .X(_2532_));
 sky130_fd_sc_hd__mux4_1 _4966_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ),
    .S0(net416),
    .S1(net406),
    .X(_2533_));
 sky130_fd_sc_hd__mux2_1 _4967_ (.A0(_2532_),
    .A1(_2533_),
    .S(net402),
    .X(_2534_));
 sky130_fd_sc_hd__mux4_1 _4968_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ),
    .S0(net418),
    .S1(net406),
    .X(_2535_));
 sky130_fd_sc_hd__mux4_1 _4969_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ),
    .S0(net418),
    .S1(net406),
    .X(_2536_));
 sky130_fd_sc_hd__mux2_1 _4970_ (.A0(_2536_),
    .A1(_2535_),
    .S(net402),
    .X(_2537_));
 sky130_fd_sc_hd__mux2_1 _4971_ (.A0(_2537_),
    .A1(_2534_),
    .S(net397),
    .X(_0051_));
 sky130_fd_sc_hd__mux4_1 _4972_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ),
    .S0(net419),
    .S1(net407),
    .X(_2538_));
 sky130_fd_sc_hd__mux4_1 _4973_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ),
    .S0(net419),
    .S1(net408),
    .X(_2539_));
 sky130_fd_sc_hd__mux2_1 _4974_ (.A0(_2538_),
    .A1(_2539_),
    .S(net401),
    .X(_2540_));
 sky130_fd_sc_hd__mux4_1 _4975_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ),
    .S0(net419),
    .S1(net408),
    .X(_2541_));
 sky130_fd_sc_hd__mux4_1 _4976_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ),
    .S0(net419),
    .S1(net408),
    .X(_2542_));
 sky130_fd_sc_hd__mux2_1 _4977_ (.A0(_2542_),
    .A1(_2541_),
    .S(net401),
    .X(_2543_));
 sky130_fd_sc_hd__mux2_1 _4978_ (.A0(_2543_),
    .A1(_2540_),
    .S(net397),
    .X(_0052_));
 sky130_fd_sc_hd__mux4_1 _4979_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ),
    .S0(net418),
    .S1(net409),
    .X(_2544_));
 sky130_fd_sc_hd__mux4_1 _4980_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ),
    .S0(net418),
    .S1(net409),
    .X(_2545_));
 sky130_fd_sc_hd__mux2_1 _4981_ (.A0(_2544_),
    .A1(_2545_),
    .S(net402),
    .X(_2546_));
 sky130_fd_sc_hd__mux4_1 _4982_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ),
    .S0(net418),
    .S1(net409),
    .X(_2547_));
 sky130_fd_sc_hd__mux4_1 _4983_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ),
    .S0(net418),
    .S1(net409),
    .X(_2548_));
 sky130_fd_sc_hd__mux2_1 _4984_ (.A0(_2548_),
    .A1(_2547_),
    .S(net402),
    .X(_2549_));
 sky130_fd_sc_hd__mux2_1 _4985_ (.A0(_2549_),
    .A1(_2546_),
    .S(net399),
    .X(_0053_));
 sky130_fd_sc_hd__mux4_1 _4986_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ),
    .S0(net417),
    .S1(net407),
    .X(_2550_));
 sky130_fd_sc_hd__mux4_1 _4987_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ),
    .S0(net417),
    .S1(net407),
    .X(_2551_));
 sky130_fd_sc_hd__mux2_1 _4988_ (.A0(_2550_),
    .A1(_2551_),
    .S(net401),
    .X(_2552_));
 sky130_fd_sc_hd__mux4_1 _4989_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ),
    .S0(net416),
    .S1(net405),
    .X(_2553_));
 sky130_fd_sc_hd__mux4_1 _4990_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ),
    .S0(net416),
    .S1(net405),
    .X(_2554_));
 sky130_fd_sc_hd__mux2_1 _4991_ (.A0(_2554_),
    .A1(_2553_),
    .S(net400),
    .X(_2555_));
 sky130_fd_sc_hd__mux2_1 _4992_ (.A0(_2555_),
    .A1(_2552_),
    .S(net397),
    .X(_0055_));
 sky130_fd_sc_hd__mux4_1 _4993_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ),
    .S0(net421),
    .S1(net411),
    .X(_2556_));
 sky130_fd_sc_hd__mux4_1 _4994_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ),
    .S0(net424),
    .S1(net411),
    .X(_2557_));
 sky130_fd_sc_hd__mux2_1 _4995_ (.A0(_2556_),
    .A1(_2557_),
    .S(net403),
    .X(_2558_));
 sky130_fd_sc_hd__mux4_1 _4996_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ),
    .S0(net420),
    .S1(net411),
    .X(_2559_));
 sky130_fd_sc_hd__mux4_1 _4997_ (.A0(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ),
    .A1(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ),
    .A2(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ),
    .A3(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ),
    .S0(net421),
    .S1(net411),
    .X(_2560_));
 sky130_fd_sc_hd__mux2_1 _4998_ (.A0(_2560_),
    .A1(_2559_),
    .S(net403),
    .X(_2561_));
 sky130_fd_sc_hd__mux2_1 _4999_ (.A0(_2561_),
    .A1(_2558_),
    .S(net397),
    .X(_0056_));
 sky130_fd_sc_hd__and2_1 _5000_ (.A(net455),
    .B(net801),
    .X(_0290_));
 sky130_fd_sc_hd__and2_1 _5001_ (.A(net455),
    .B(net743),
    .X(_0291_));
 sky130_fd_sc_hd__and2_4 _5002_ (.A(net439),
    .B(net171),
    .X(_2562_));
 sky130_fd_sc_hd__mux2_1 _5003_ (.A0(net2122),
    .A1(net925),
    .S(net239),
    .X(_2563_));
 sky130_fd_sc_hd__or3b_1 _5004_ (.A(net468),
    .B(_2563_),
    .C_N(net2117),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _5005_ (.A(net1013),
    .B(net226),
    .X(_2564_));
 sky130_fd_sc_hd__o211a_1 _5006_ (.A1(net2024),
    .A2(net238),
    .B1(net165),
    .C1(_2564_),
    .X(_0323_));
 sky130_fd_sc_hd__or2_1 _5007_ (.A(net839),
    .B(net221),
    .X(_2565_));
 sky130_fd_sc_hd__o211a_1 _5008_ (.A1(net2068),
    .A2(net237),
    .B1(net163),
    .C1(_2565_),
    .X(_0324_));
 sky130_fd_sc_hd__or2_1 _5009_ (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[5] ),
    .B(net221),
    .X(_2566_));
 sky130_fd_sc_hd__o211a_1 _5010_ (.A1(net837),
    .A2(net236),
    .B1(net163),
    .C1(_2566_),
    .X(_0325_));
 sky130_fd_sc_hd__or2_1 _5011_ (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ),
    .B(net227),
    .X(_2567_));
 sky130_fd_sc_hd__o211a_1 _5012_ (.A1(net817),
    .A2(net239),
    .B1(net165),
    .C1(_2567_),
    .X(_0326_));
 sky130_fd_sc_hd__or2_1 _5013_ (.A(net883),
    .B(net225),
    .X(_2568_));
 sky130_fd_sc_hd__o211a_1 _5014_ (.A1(net2065),
    .A2(net238),
    .B1(net165),
    .C1(_2568_),
    .X(_0327_));
 sky130_fd_sc_hd__or2_1 _5015_ (.A(net897),
    .B(net227),
    .X(_2569_));
 sky130_fd_sc_hd__o211a_1 _5016_ (.A1(net1893),
    .A2(net238),
    .B1(net165),
    .C1(_2569_),
    .X(_0328_));
 sky130_fd_sc_hd__or2_1 _5017_ (.A(net969),
    .B(net231),
    .X(_2570_));
 sky130_fd_sc_hd__o211a_1 _5018_ (.A1(net1998),
    .A2(net240),
    .B1(net164),
    .C1(_2570_),
    .X(_0329_));
 sky130_fd_sc_hd__or2_1 _5019_ (.A(net877),
    .B(net230),
    .X(_2571_));
 sky130_fd_sc_hd__o211a_1 _5020_ (.A1(net1994),
    .A2(net240),
    .B1(net164),
    .C1(_2571_),
    .X(_0330_));
 sky130_fd_sc_hd__or2_1 _5021_ (.A(net849),
    .B(net229),
    .X(_2572_));
 sky130_fd_sc_hd__o211a_1 _5022_ (.A1(net2022),
    .A2(net241),
    .B1(net164),
    .C1(_2572_),
    .X(_0331_));
 sky130_fd_sc_hd__or2_1 _5023_ (.A(net931),
    .B(net231),
    .X(_2573_));
 sky130_fd_sc_hd__o211a_1 _5024_ (.A1(net2003),
    .A2(net240),
    .B1(net166),
    .C1(_2573_),
    .X(_0332_));
 sky130_fd_sc_hd__or2_1 _5025_ (.A(net943),
    .B(net230),
    .X(_2574_));
 sky130_fd_sc_hd__o211a_1 _5026_ (.A1(net1792),
    .A2(net240),
    .B1(net166),
    .C1(_2574_),
    .X(_0333_));
 sky130_fd_sc_hd__or2_1 _5027_ (.A(net973),
    .B(net230),
    .X(_2575_));
 sky130_fd_sc_hd__o211a_1 _5028_ (.A1(net1242),
    .A2(net240),
    .B1(net166),
    .C1(_2575_),
    .X(_0334_));
 sky130_fd_sc_hd__or2_1 _5029_ (.A(net1152),
    .B(net214),
    .X(_2576_));
 sky130_fd_sc_hd__o211a_1 _5030_ (.A1(net2036),
    .A2(net233),
    .B1(net161),
    .C1(_2576_),
    .X(_0335_));
 sky130_fd_sc_hd__or2_1 _5031_ (.A(net921),
    .B(net214),
    .X(_2577_));
 sky130_fd_sc_hd__o211a_1 _5032_ (.A1(net1997),
    .A2(net233),
    .B1(net161),
    .C1(_2577_),
    .X(_0336_));
 sky130_fd_sc_hd__or2_1 _5033_ (.A(net951),
    .B(net215),
    .X(_2578_));
 sky130_fd_sc_hd__o211a_1 _5034_ (.A1(net1984),
    .A2(net233),
    .B1(net161),
    .C1(_2578_),
    .X(_0337_));
 sky130_fd_sc_hd__or2_1 _5035_ (.A(net985),
    .B(net217),
    .X(_2579_));
 sky130_fd_sc_hd__o211a_1 _5036_ (.A1(net1987),
    .A2(net235),
    .B1(net162),
    .C1(_2579_),
    .X(_0338_));
 sky130_fd_sc_hd__or2_1 _5037_ (.A(net1322),
    .B(net216),
    .X(_2580_));
 sky130_fd_sc_hd__o211a_1 _5038_ (.A1(net1784),
    .A2(net234),
    .B1(net161),
    .C1(_2580_),
    .X(_0339_));
 sky130_fd_sc_hd__or2_1 _5039_ (.A(net809),
    .B(net218),
    .X(_2581_));
 sky130_fd_sc_hd__o211a_1 _5040_ (.A1(net2019),
    .A2(net235),
    .B1(net162),
    .C1(_2581_),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _5041_ (.A(net783),
    .B(net219),
    .X(_2582_));
 sky130_fd_sc_hd__o211a_1 _5042_ (.A1(net1969),
    .A2(net234),
    .B1(net161),
    .C1(_2582_),
    .X(_0341_));
 sky130_fd_sc_hd__or2_1 _5043_ (.A(net803),
    .B(net214),
    .X(_2583_));
 sky130_fd_sc_hd__o211a_1 _5044_ (.A1(net1820),
    .A2(net233),
    .B1(net161),
    .C1(_2583_),
    .X(_0342_));
 sky130_fd_sc_hd__or2_1 _5045_ (.A(net821),
    .B(net215),
    .X(_2584_));
 sky130_fd_sc_hd__o211a_1 _5046_ (.A1(net2038),
    .A2(net233),
    .B1(net161),
    .C1(_2584_),
    .X(_0343_));
 sky130_fd_sc_hd__or2_1 _5047_ (.A(net901),
    .B(net218),
    .X(_2585_));
 sky130_fd_sc_hd__o211a_1 _5048_ (.A1(net2000),
    .A2(net235),
    .B1(net161),
    .C1(_2585_),
    .X(_0344_));
 sky130_fd_sc_hd__or2_1 _5049_ (.A(net703),
    .B(net217),
    .X(_2586_));
 sky130_fd_sc_hd__o211a_1 _5050_ (.A1(net2017),
    .A2(net235),
    .B1(net162),
    .C1(_2586_),
    .X(_0345_));
 sky130_fd_sc_hd__or2_1 _5051_ (.A(net893),
    .B(net217),
    .X(_2587_));
 sky130_fd_sc_hd__o211a_1 _5052_ (.A1(net1993),
    .A2(net235),
    .B1(net161),
    .C1(_2587_),
    .X(_0346_));
 sky130_fd_sc_hd__or2_1 _5053_ (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[27] ),
    .B(net220),
    .X(_2588_));
 sky130_fd_sc_hd__o211a_1 _5054_ (.A1(net871),
    .A2(net236),
    .B1(net163),
    .C1(_2588_),
    .X(_0347_));
 sky130_fd_sc_hd__or2_1 _5055_ (.A(net913),
    .B(net220),
    .X(_2589_));
 sky130_fd_sc_hd__o211a_1 _5056_ (.A1(net2011),
    .A2(net236),
    .B1(net163),
    .C1(_2589_),
    .X(_0348_));
 sky130_fd_sc_hd__or2_1 _5057_ (.A(net955),
    .B(net222),
    .X(_2590_));
 sky130_fd_sc_hd__o211a_1 _5058_ (.A1(net2008),
    .A2(net236),
    .B1(net163),
    .C1(_2590_),
    .X(_0349_));
 sky130_fd_sc_hd__or2_1 _5059_ (.A(net989),
    .B(net222),
    .X(_2591_));
 sky130_fd_sc_hd__o211a_1 _5060_ (.A1(net1983),
    .A2(net236),
    .B1(net163),
    .C1(_2591_),
    .X(_0350_));
 sky130_fd_sc_hd__or2_1 _5061_ (.A(net941),
    .B(net221),
    .X(_2592_));
 sky130_fd_sc_hd__o211a_1 _5062_ (.A1(net1990),
    .A2(net237),
    .B1(net163),
    .C1(_2592_),
    .X(_0351_));
 sky130_fd_sc_hd__or2_1 _5063_ (.A(net2254),
    .B(net231),
    .X(_2593_));
 sky130_fd_sc_hd__o211a_1 _5064_ (.A1(net21),
    .A2(net240),
    .B1(net164),
    .C1(_2593_),
    .X(_0352_));
 sky130_fd_sc_hd__or2_1 _5065_ (.A(net2210),
    .B(net218),
    .X(_2594_));
 sky130_fd_sc_hd__o211a_1 _5066_ (.A1(net24),
    .A2(net235),
    .B1(net162),
    .C1(_2594_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _5067_ (.A0(net25),
    .A1(net2258),
    .S(net235),
    .X(_2595_));
 sky130_fd_sc_hd__or3b_1 _5068_ (.A(net463),
    .B(_2595_),
    .C_N(net171),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _5069_ (.A0(net26),
    .A1(net2170),
    .S(net236),
    .X(_2596_));
 sky130_fd_sc_hd__or3b_1 _5070_ (.A(net464),
    .B(_2596_),
    .C_N(net172),
    .X(_0355_));
 sky130_fd_sc_hd__or2_1 _5071_ (.A(net1988),
    .B(net225),
    .X(_2597_));
 sky130_fd_sc_hd__o211a_1 _5072_ (.A1(net27),
    .A2(net238),
    .B1(net165),
    .C1(_2597_),
    .X(_0356_));
 sky130_fd_sc_hd__nand2_1 _5073_ (.A(_1404_),
    .B(net239),
    .Y(_2598_));
 sky130_fd_sc_hd__o211a_1 _5074_ (.A1(net28),
    .A2(net239),
    .B1(net165),
    .C1(_2598_),
    .X(_0357_));
 sky130_fd_sc_hd__or2_1 _5075_ (.A(net1991),
    .B(net224),
    .X(_2599_));
 sky130_fd_sc_hd__o211a_1 _5076_ (.A1(net29),
    .A2(net242),
    .B1(net166),
    .C1(_2599_),
    .X(_0358_));
 sky130_fd_sc_hd__or2_1 _5077_ (.A(net2121),
    .B(net229),
    .X(_2600_));
 sky130_fd_sc_hd__o211a_1 _5078_ (.A1(net30),
    .A2(net241),
    .B1(net164),
    .C1(_2600_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _5079_ (.A(net2118),
    .B(net229),
    .X(_2601_));
 sky130_fd_sc_hd__o211a_1 _5080_ (.A1(net1),
    .A2(net241),
    .B1(net164),
    .C1(_2601_),
    .X(_0360_));
 sky130_fd_sc_hd__or2_1 _5081_ (.A(net2198),
    .B(net227),
    .X(_2602_));
 sky130_fd_sc_hd__o211a_1 _5082_ (.A1(net2),
    .A2(net238),
    .B1(net165),
    .C1(_2602_),
    .X(_0361_));
 sky130_fd_sc_hd__or2_1 _5083_ (.A(net2127),
    .B(net229),
    .X(_2603_));
 sky130_fd_sc_hd__o211a_1 _5084_ (.A1(net3),
    .A2(net241),
    .B1(net164),
    .C1(_2603_),
    .X(_0362_));
 sky130_fd_sc_hd__nand2_1 _5085_ (.A(_1403_),
    .B(net239),
    .Y(_2604_));
 sky130_fd_sc_hd__o211a_1 _5086_ (.A1(net4),
    .A2(net239),
    .B1(net165),
    .C1(_2604_),
    .X(_0363_));
 sky130_fd_sc_hd__or2_1 _5087_ (.A(net2145),
    .B(net231),
    .X(_2605_));
 sky130_fd_sc_hd__o211a_1 _5088_ (.A1(net5),
    .A2(net240),
    .B1(net164),
    .C1(_2605_),
    .X(_0364_));
 sky130_fd_sc_hd__or2_1 _5089_ (.A(net415),
    .B(net213),
    .X(_2606_));
 sky130_fd_sc_hd__o211a_1 _5090_ (.A1(net6),
    .A2(net242),
    .B1(_2562_),
    .C1(_2606_),
    .X(_0365_));
 sky130_fd_sc_hd__or2_1 _5091_ (.A(net409),
    .B(net218),
    .X(_2607_));
 sky130_fd_sc_hd__o211a_1 _5092_ (.A1(net7),
    .A2(net235),
    .B1(net162),
    .C1(_2607_),
    .X(_0366_));
 sky130_fd_sc_hd__or2_1 _5093_ (.A(net404),
    .B(net229),
    .X(_2608_));
 sky130_fd_sc_hd__o211a_1 _5094_ (.A1(net8),
    .A2(net241),
    .B1(net164),
    .C1(_2608_),
    .X(_0367_));
 sky130_fd_sc_hd__or2_1 _5095_ (.A(net399),
    .B(net217),
    .X(_2609_));
 sky130_fd_sc_hd__o211a_1 _5096_ (.A1(net9),
    .A2(net235),
    .B1(net162),
    .C1(_2609_),
    .X(_0368_));
 sky130_fd_sc_hd__or2_1 _5097_ (.A(net694),
    .B(net221),
    .X(_2610_));
 sky130_fd_sc_hd__o211a_1 _5098_ (.A1(net10),
    .A2(net238),
    .B1(net165),
    .C1(_2610_),
    .X(_0369_));
 sky130_fd_sc_hd__nand2_1 _5099_ (.A(_1402_),
    .B(net242),
    .Y(_2611_));
 sky130_fd_sc_hd__o211a_1 _5100_ (.A1(net11),
    .A2(net242),
    .B1(_2562_),
    .C1(_2611_),
    .X(_0370_));
 sky130_fd_sc_hd__or2_1 _5101_ (.A(net385),
    .B(net224),
    .X(_2612_));
 sky130_fd_sc_hd__o211a_1 _5102_ (.A1(net12),
    .A2(net242),
    .B1(net166),
    .C1(_2612_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _5103_ (.A(net370),
    .B(net213),
    .X(_2613_));
 sky130_fd_sc_hd__o211a_1 _5104_ (.A1(net13),
    .A2(net242),
    .B1(_2562_),
    .C1(_2613_),
    .X(_0372_));
 sky130_fd_sc_hd__or2_1 _5105_ (.A(net369),
    .B(net223),
    .X(_2614_));
 sky130_fd_sc_hd__o211a_1 _5106_ (.A1(net14),
    .A2(net242),
    .B1(net166),
    .C1(_2614_),
    .X(_0373_));
 sky130_fd_sc_hd__or2_1 _5107_ (.A(net2109),
    .B(net213),
    .X(_2615_));
 sky130_fd_sc_hd__o211a_1 _5108_ (.A1(net15),
    .A2(net242),
    .B1(_2562_),
    .C1(_2615_),
    .X(_0374_));
 sky130_fd_sc_hd__or2_1 _5109_ (.A(net2083),
    .B(net221),
    .X(_2616_));
 sky130_fd_sc_hd__o211a_1 _5110_ (.A1(net16),
    .A2(net236),
    .B1(net163),
    .C1(_2616_),
    .X(_0375_));
 sky130_fd_sc_hd__or2_1 _5111_ (.A(net2188),
    .B(net224),
    .X(_2617_));
 sky130_fd_sc_hd__o211a_1 _5112_ (.A1(net17),
    .A2(net242),
    .B1(net166),
    .C1(_2617_),
    .X(_0376_));
 sky130_fd_sc_hd__or2_1 _5113_ (.A(net1878),
    .B(net229),
    .X(_2618_));
 sky130_fd_sc_hd__o211a_1 _5114_ (.A1(net18),
    .A2(net241),
    .B1(net164),
    .C1(_2618_),
    .X(_0377_));
 sky130_fd_sc_hd__or2_1 _5115_ (.A(net2175),
    .B(net223),
    .X(_2619_));
 sky130_fd_sc_hd__o211a_1 _5116_ (.A1(net19),
    .A2(net242),
    .B1(net166),
    .C1(_2619_),
    .X(_0378_));
 sky130_fd_sc_hd__or2_1 _5117_ (.A(net1971),
    .B(net218),
    .X(_2620_));
 sky130_fd_sc_hd__o211a_1 _5118_ (.A1(net20),
    .A2(net235),
    .B1(net162),
    .C1(_2620_),
    .X(_0379_));
 sky130_fd_sc_hd__or2_1 _5119_ (.A(net2048),
    .B(net228),
    .X(_2621_));
 sky130_fd_sc_hd__o211a_1 _5120_ (.A1(net22),
    .A2(net241),
    .B1(net164),
    .C1(_2621_),
    .X(_0380_));
 sky130_fd_sc_hd__or2_1 _5121_ (.A(net2090),
    .B(net229),
    .X(_2622_));
 sky130_fd_sc_hd__o211a_1 _5122_ (.A1(net23),
    .A2(net241),
    .B1(net164),
    .C1(_2622_),
    .X(_0381_));
 sky130_fd_sc_hd__or2_1 _5123_ (.A(net887),
    .B(net225),
    .X(_2623_));
 sky130_fd_sc_hd__o211a_1 _5124_ (.A1(net2057),
    .A2(net238),
    .B1(net165),
    .C1(_2623_),
    .X(_0382_));
 sky130_fd_sc_hd__or2_1 _5125_ (.A(net873),
    .B(net226),
    .X(_2624_));
 sky130_fd_sc_hd__o211a_1 _5126_ (.A1(net2051),
    .A2(net238),
    .B1(net165),
    .C1(_2624_),
    .X(_0383_));
 sky130_fd_sc_hd__or2_1 _5127_ (.A(net819),
    .B(net221),
    .X(_2625_));
 sky130_fd_sc_hd__o211a_1 _5128_ (.A1(net2072),
    .A2(net237),
    .B1(net163),
    .C1(_2625_),
    .X(_0384_));
 sky130_fd_sc_hd__or2_1 _5129_ (.A(net827),
    .B(net225),
    .X(_2626_));
 sky130_fd_sc_hd__o211a_1 _5130_ (.A1(net2058),
    .A2(net238),
    .B1(net165),
    .C1(_2626_),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _5131_ (.A(net1130),
    .B(net225),
    .X(_2627_));
 sky130_fd_sc_hd__o211a_1 _5132_ (.A1(net2103),
    .A2(net238),
    .B1(net165),
    .C1(_2627_),
    .X(_0386_));
 sky130_fd_sc_hd__or2_1 _5133_ (.A(net875),
    .B(net225),
    .X(_2628_));
 sky130_fd_sc_hd__o211a_1 _5134_ (.A1(net2044),
    .A2(net238),
    .B1(net165),
    .C1(_2628_),
    .X(_0387_));
 sky130_fd_sc_hd__or2_1 _5135_ (.A(net853),
    .B(net227),
    .X(_2629_));
 sky130_fd_sc_hd__o211a_1 _5136_ (.A1(net2064),
    .A2(net239),
    .B1(net165),
    .C1(_2629_),
    .X(_0388_));
 sky130_fd_sc_hd__or2_1 _5137_ (.A(net823),
    .B(net230),
    .X(_2630_));
 sky130_fd_sc_hd__o211a_1 _5138_ (.A1(net2073),
    .A2(net240),
    .B1(net164),
    .C1(_2630_),
    .X(_0389_));
 sky130_fd_sc_hd__or2_1 _5139_ (.A(net961),
    .B(net227),
    .X(_2631_));
 sky130_fd_sc_hd__o211a_1 _5140_ (.A1(net2074),
    .A2(net238),
    .B1(net165),
    .C1(_2631_),
    .X(_0390_));
 sky130_fd_sc_hd__or2_1 _5141_ (.A(net987),
    .B(net228),
    .X(_2632_));
 sky130_fd_sc_hd__o211a_1 _5142_ (.A1(net2081),
    .A2(net241),
    .B1(net164),
    .C1(_2632_),
    .X(_0391_));
 sky130_fd_sc_hd__or2_1 _5143_ (.A(net937),
    .B(net231),
    .X(_2633_));
 sky130_fd_sc_hd__o211a_1 _5144_ (.A1(net2079),
    .A2(net241),
    .B1(net164),
    .C1(_2633_),
    .X(_0392_));
 sky130_fd_sc_hd__or2_1 _5145_ (.A(net899),
    .B(net230),
    .X(_2634_));
 sky130_fd_sc_hd__o211a_1 _5146_ (.A1(net2046),
    .A2(net240),
    .B1(net164),
    .C1(_2634_),
    .X(_0393_));
 sky130_fd_sc_hd__or2_1 _5147_ (.A(net967),
    .B(net231),
    .X(_2635_));
 sky130_fd_sc_hd__o211a_1 _5148_ (.A1(net2088),
    .A2(net240),
    .B1(net166),
    .C1(_2635_),
    .X(_0394_));
 sky130_fd_sc_hd__or2_1 _5149_ (.A(net995),
    .B(net214),
    .X(_2636_));
 sky130_fd_sc_hd__o211a_1 _5150_ (.A1(net2108),
    .A2(net233),
    .B1(net161),
    .C1(_2636_),
    .X(_0395_));
 sky130_fd_sc_hd__or2_1 _5151_ (.A(net979),
    .B(net216),
    .X(_2637_));
 sky130_fd_sc_hd__o211a_1 _5152_ (.A1(net2089),
    .A2(net234),
    .B1(net161),
    .C1(_2637_),
    .X(_0396_));
 sky130_fd_sc_hd__or2_1 _5153_ (.A(net993),
    .B(net216),
    .X(_2638_));
 sky130_fd_sc_hd__o211a_1 _5154_ (.A1(net2086),
    .A2(net234),
    .B1(net161),
    .C1(_2638_),
    .X(_0397_));
 sky130_fd_sc_hd__or2_1 _5155_ (.A(net813),
    .B(net216),
    .X(_2639_));
 sky130_fd_sc_hd__o211a_1 _5156_ (.A1(net2075),
    .A2(net233),
    .B1(net161),
    .C1(_2639_),
    .X(_0398_));
 sky130_fd_sc_hd__or2_1 _5157_ (.A(net1104),
    .B(net217),
    .X(_2640_));
 sky130_fd_sc_hd__o211a_1 _5158_ (.A1(net2078),
    .A2(net236),
    .B1(_2562_),
    .C1(_2640_),
    .X(_0399_));
 sky130_fd_sc_hd__or2_1 _5159_ (.A(net915),
    .B(net214),
    .X(_2641_));
 sky130_fd_sc_hd__o211a_1 _5160_ (.A1(net2059),
    .A2(net233),
    .B1(net161),
    .C1(_2641_),
    .X(_0400_));
 sky130_fd_sc_hd__or2_1 _5161_ (.A(net648),
    .B(net217),
    .X(_2642_));
 sky130_fd_sc_hd__o211a_1 _5162_ (.A1(net2047),
    .A2(net235),
    .B1(net162),
    .C1(_2642_),
    .X(_0401_));
 sky130_fd_sc_hd__or2_1 _5163_ (.A(net855),
    .B(net216),
    .X(_2643_));
 sky130_fd_sc_hd__o211a_1 _5164_ (.A1(net2034),
    .A2(net233),
    .B1(net161),
    .C1(_2643_),
    .X(_0402_));
 sky130_fd_sc_hd__or2_1 _5165_ (.A(net929),
    .B(net214),
    .X(_2644_));
 sky130_fd_sc_hd__o211a_1 _5166_ (.A1(net2069),
    .A2(net233),
    .B1(net161),
    .C1(_2644_),
    .X(_0403_));
 sky130_fd_sc_hd__or2_1 _5167_ (.A(net911),
    .B(net217),
    .X(_2645_));
 sky130_fd_sc_hd__o211a_1 _5168_ (.A1(net2067),
    .A2(net235),
    .B1(net162),
    .C1(_2645_),
    .X(_0404_));
 sky130_fd_sc_hd__or2_1 _5169_ (.A(net907),
    .B(net218),
    .X(_2646_));
 sky130_fd_sc_hd__o211a_1 _5170_ (.A1(net2082),
    .A2(net235),
    .B1(net162),
    .C1(_2646_),
    .X(_0405_));
 sky130_fd_sc_hd__or2_1 _5171_ (.A(net670),
    .B(net217),
    .X(_2647_));
 sky130_fd_sc_hd__o211a_1 _5172_ (.A1(net2080),
    .A2(net235),
    .B1(net162),
    .C1(_2647_),
    .X(_0406_));
 sky130_fd_sc_hd__or2_1 _5173_ (.A(net668),
    .B(net220),
    .X(_2648_));
 sky130_fd_sc_hd__o211a_1 _5174_ (.A1(net2097),
    .A2(net236),
    .B1(net163),
    .C1(_2648_),
    .X(_0407_));
 sky130_fd_sc_hd__or2_1 _5175_ (.A(net672),
    .B(net220),
    .X(_2649_));
 sky130_fd_sc_hd__o211a_1 _5176_ (.A1(net2096),
    .A2(net236),
    .B1(net163),
    .C1(_2649_),
    .X(_0408_));
 sky130_fd_sc_hd__or2_1 _5177_ (.A(net1098),
    .B(net220),
    .X(_2650_));
 sky130_fd_sc_hd__o211a_1 _5178_ (.A1(net2093),
    .A2(net236),
    .B1(net163),
    .C1(_2650_),
    .X(_0409_));
 sky130_fd_sc_hd__or2_1 _5179_ (.A(net933),
    .B(net222),
    .X(_2651_));
 sky130_fd_sc_hd__o211a_1 _5180_ (.A1(net2070),
    .A2(net237),
    .B1(net163),
    .C1(_2651_),
    .X(_0410_));
 sky130_fd_sc_hd__or2_1 _5181_ (.A(net1310),
    .B(net222),
    .X(_2652_));
 sky130_fd_sc_hd__o211a_1 _5182_ (.A1(net2098),
    .A2(net237),
    .B1(net163),
    .C1(_2652_),
    .X(_0411_));
 sky130_fd_sc_hd__and2_1 _5183_ (.A(net453),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ),
    .X(_2653_));
 sky130_fd_sc_hd__or3b_4 _5184_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(_1408_),
    .C_N(_2653_),
    .X(_2654_));
 sky130_fd_sc_hd__nand2_4 _5185_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .Y(_2655_));
 sky130_fd_sc_hd__nor2_2 _5186_ (.A(_2654_),
    .B(_2655_),
    .Y(_2656_));
 sky130_fd_sc_hd__or2_1 _5187_ (.A(_2654_),
    .B(_2655_),
    .X(_2657_));
 sky130_fd_sc_hd__nor2_1 _5188_ (.A(net466),
    .B(net315),
    .Y(_2658_));
 sky130_fd_sc_hd__nand2_1 _5189_ (.A(net450),
    .B(_2657_),
    .Y(_2659_));
 sky130_fd_sc_hd__a22o_1 _5190_ (.A1(net356),
    .A2(net316),
    .B1(net266),
    .B2(net1148),
    .X(_0412_));
 sky130_fd_sc_hd__o22a_1 _5191_ (.A1(_1689_),
    .A2(_2657_),
    .B1(_2659_),
    .B2(net949),
    .X(_0413_));
 sky130_fd_sc_hd__o22a_1 _5192_ (.A1(net329),
    .A2(_2657_),
    .B1(_2659_),
    .B2(net891),
    .X(_0414_));
 sky130_fd_sc_hd__o22a_1 _5193_ (.A1(net330),
    .A2(_2657_),
    .B1(_2659_),
    .B2(net889),
    .X(_0415_));
 sky130_fd_sc_hd__a22o_1 _5194_ (.A1(net327),
    .A2(net315),
    .B1(net265),
    .B2(net1688),
    .X(_0416_));
 sky130_fd_sc_hd__a22o_1 _5195_ (.A1(net325),
    .A2(net316),
    .B1(net266),
    .B2(net1078),
    .X(_0417_));
 sky130_fd_sc_hd__a22o_1 _5196_ (.A1(net328),
    .A2(net316),
    .B1(net266),
    .B2(net1272),
    .X(_0418_));
 sky130_fd_sc_hd__a22o_1 _5197_ (.A1(net326),
    .A2(net315),
    .B1(net265),
    .B2(net1638),
    .X(_0419_));
 sky130_fd_sc_hd__a22o_1 _5198_ (.A1(net323),
    .A2(net316),
    .B1(net266),
    .B2(net1646),
    .X(_0420_));
 sky130_fd_sc_hd__a22o_1 _5199_ (.A1(net321),
    .A2(net316),
    .B1(net266),
    .B2(net1426),
    .X(_0421_));
 sky130_fd_sc_hd__a22o_1 _5200_ (.A1(net324),
    .A2(net316),
    .B1(net266),
    .B2(net1462),
    .X(_0422_));
 sky130_fd_sc_hd__a22o_1 _5201_ (.A1(net322),
    .A2(net315),
    .B1(net265),
    .B2(net1226),
    .X(_0423_));
 sky130_fd_sc_hd__a22o_1 _5202_ (.A1(net319),
    .A2(net316),
    .B1(net266),
    .B2(net1274),
    .X(_0424_));
 sky130_fd_sc_hd__a22o_1 _5203_ (.A1(_1832_),
    .A2(net316),
    .B1(net266),
    .B2(net1536),
    .X(_0425_));
 sky130_fd_sc_hd__a22o_1 _5204_ (.A1(net320),
    .A2(net316),
    .B1(net266),
    .B2(net1356),
    .X(_0426_));
 sky130_fd_sc_hd__a22o_1 _5205_ (.A1(net318),
    .A2(net315),
    .B1(net265),
    .B2(net1110),
    .X(_0427_));
 sky130_fd_sc_hd__a22o_1 _5206_ (.A1(net341),
    .A2(net316),
    .B1(net265),
    .B2(net1052),
    .X(_0428_));
 sky130_fd_sc_hd__a22o_1 _5207_ (.A1(net340),
    .A2(net316),
    .B1(net266),
    .B2(net1414),
    .X(_0429_));
 sky130_fd_sc_hd__a22o_1 _5208_ (.A1(net339),
    .A2(net315),
    .B1(net265),
    .B2(net1438),
    .X(_0430_));
 sky130_fd_sc_hd__a22o_1 _5209_ (.A1(net338),
    .A2(net315),
    .B1(net265),
    .B2(net1602),
    .X(_0431_));
 sky130_fd_sc_hd__a22o_1 _5210_ (.A1(net333),
    .A2(net315),
    .B1(net265),
    .B2(net1278),
    .X(_0432_));
 sky130_fd_sc_hd__a22o_1 _5211_ (.A1(net331),
    .A2(net316),
    .B1(net266),
    .B2(net1244),
    .X(_0433_));
 sky130_fd_sc_hd__a22o_1 _5212_ (.A1(net334),
    .A2(net315),
    .B1(net265),
    .B2(net1454),
    .X(_0434_));
 sky130_fd_sc_hd__a22o_1 _5213_ (.A1(net332),
    .A2(net315),
    .B1(net265),
    .B2(net1214),
    .X(_0435_));
 sky130_fd_sc_hd__a22o_1 _5214_ (.A1(net343),
    .A2(net315),
    .B1(net265),
    .B2(net1208),
    .X(_0436_));
 sky130_fd_sc_hd__a22o_1 _5215_ (.A1(net348),
    .A2(net316),
    .B1(net266),
    .B2(net1364),
    .X(_0437_));
 sky130_fd_sc_hd__a22o_1 _5216_ (.A1(net344),
    .A2(net315),
    .B1(net265),
    .B2(net1106),
    .X(_0438_));
 sky130_fd_sc_hd__a22o_1 _5217_ (.A1(net342),
    .A2(net315),
    .B1(net265),
    .B2(net1072),
    .X(_0439_));
 sky130_fd_sc_hd__a22o_1 _5218_ (.A1(net336),
    .A2(net315),
    .B1(net265),
    .B2(net1560),
    .X(_0440_));
 sky130_fd_sc_hd__a22o_1 _5219_ (.A1(net335),
    .A2(net315),
    .B1(net265),
    .B2(net1622),
    .X(_0441_));
 sky130_fd_sc_hd__a22o_1 _5220_ (.A1(net337),
    .A2(net315),
    .B1(net265),
    .B2(net1340),
    .X(_0442_));
 sky130_fd_sc_hd__a22o_1 _5221_ (.A1(net357),
    .A2(net316),
    .B1(net266),
    .B2(net1522),
    .X(_0443_));
 sky130_fd_sc_hd__or3b_4 _5222_ (.A(_1407_),
    .B(_1408_),
    .C_N(_2653_),
    .X(_2660_));
 sky130_fd_sc_hd__nand2_4 _5223_ (.A(_1409_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .Y(_2661_));
 sky130_fd_sc_hd__nor2_1 _5224_ (.A(_2660_),
    .B(_2661_),
    .Y(_2662_));
 sky130_fd_sc_hd__or2_1 _5225_ (.A(_2660_),
    .B(_2661_),
    .X(_2663_));
 sky130_fd_sc_hd__nor2_2 _5226_ (.A(net461),
    .B(net314),
    .Y(_2664_));
 sky130_fd_sc_hd__nand2_1 _5227_ (.A(net449),
    .B(_2663_),
    .Y(_2665_));
 sky130_fd_sc_hd__o22a_1 _5228_ (.A1(net356),
    .A2(_2663_),
    .B1(_2665_),
    .B2(net939),
    .X(_0444_));
 sky130_fd_sc_hd__o22a_1 _5229_ (.A1(_1689_),
    .A2(_2663_),
    .B1(_2665_),
    .B2(net963),
    .X(_0445_));
 sky130_fd_sc_hd__a22o_1 _5230_ (.A1(net329),
    .A2(net314),
    .B1(net264),
    .B2(net1380),
    .X(_0446_));
 sky130_fd_sc_hd__o22a_1 _5231_ (.A1(net330),
    .A2(_2663_),
    .B1(_2665_),
    .B2(net859),
    .X(_0447_));
 sky130_fd_sc_hd__a22o_1 _5232_ (.A1(net327),
    .A2(net313),
    .B1(net263),
    .B2(net1464),
    .X(_0448_));
 sky130_fd_sc_hd__a22o_1 _5233_ (.A1(net325),
    .A2(net314),
    .B1(net264),
    .B2(net1358),
    .X(_0449_));
 sky130_fd_sc_hd__a22o_1 _5234_ (.A1(net328),
    .A2(net314),
    .B1(net264),
    .B2(net1406),
    .X(_0450_));
 sky130_fd_sc_hd__a22o_1 _5235_ (.A1(net326),
    .A2(net313),
    .B1(net263),
    .B2(net1594),
    .X(_0451_));
 sky130_fd_sc_hd__a22o_1 _5236_ (.A1(net323),
    .A2(net314),
    .B1(net264),
    .B2(net1478),
    .X(_0452_));
 sky130_fd_sc_hd__a22o_1 _5237_ (.A1(net321),
    .A2(net314),
    .B1(net264),
    .B2(net1150),
    .X(_0453_));
 sky130_fd_sc_hd__a22o_1 _5238_ (.A1(net324),
    .A2(net314),
    .B1(net264),
    .B2(net1122),
    .X(_0454_));
 sky130_fd_sc_hd__a22o_1 _5239_ (.A1(net322),
    .A2(net313),
    .B1(net263),
    .B2(net1254),
    .X(_0455_));
 sky130_fd_sc_hd__a22o_1 _5240_ (.A1(net319),
    .A2(net314),
    .B1(net264),
    .B2(net1200),
    .X(_0456_));
 sky130_fd_sc_hd__a22o_1 _5241_ (.A1(net317),
    .A2(net314),
    .B1(net264),
    .B2(net1712),
    .X(_0457_));
 sky130_fd_sc_hd__a22o_1 _5242_ (.A1(net320),
    .A2(net314),
    .B1(net264),
    .B2(net1094),
    .X(_0458_));
 sky130_fd_sc_hd__a22o_1 _5243_ (.A1(net318),
    .A2(net313),
    .B1(net263),
    .B2(net1212),
    .X(_0459_));
 sky130_fd_sc_hd__a22o_1 _5244_ (.A1(net341),
    .A2(net313),
    .B1(net263),
    .B2(net1024),
    .X(_0460_));
 sky130_fd_sc_hd__a22o_1 _5245_ (.A1(net340),
    .A2(net314),
    .B1(net264),
    .B2(net1532),
    .X(_0461_));
 sky130_fd_sc_hd__a22o_1 _5246_ (.A1(net339),
    .A2(net313),
    .B1(net263),
    .B2(net1086),
    .X(_0462_));
 sky130_fd_sc_hd__a22o_1 _5247_ (.A1(net338),
    .A2(net313),
    .B1(net263),
    .B2(net1580),
    .X(_0463_));
 sky130_fd_sc_hd__a22o_1 _5248_ (.A1(net333),
    .A2(net313),
    .B1(net263),
    .B2(net999),
    .X(_0464_));
 sky130_fd_sc_hd__a22o_1 _5249_ (.A1(net331),
    .A2(net314),
    .B1(net264),
    .B2(net1034),
    .X(_0465_));
 sky130_fd_sc_hd__a22o_1 _5250_ (.A1(net334),
    .A2(net313),
    .B1(net263),
    .B2(net1282),
    .X(_0466_));
 sky130_fd_sc_hd__a22o_1 _5251_ (.A1(net332),
    .A2(net313),
    .B1(net263),
    .B2(net1140),
    .X(_0467_));
 sky130_fd_sc_hd__a22o_1 _5252_ (.A1(net343),
    .A2(net313),
    .B1(net263),
    .B2(net1054),
    .X(_0468_));
 sky130_fd_sc_hd__a22o_1 _5253_ (.A1(net348),
    .A2(net314),
    .B1(net264),
    .B2(net981),
    .X(_0469_));
 sky130_fd_sc_hd__a22o_1 _5254_ (.A1(net344),
    .A2(net313),
    .B1(net263),
    .B2(net1154),
    .X(_0470_));
 sky130_fd_sc_hd__a22o_1 _5255_ (.A1(net342),
    .A2(net313),
    .B1(net263),
    .B2(net1058),
    .X(_0471_));
 sky130_fd_sc_hd__a22o_1 _5256_ (.A1(net336),
    .A2(net313),
    .B1(net263),
    .B2(net1306),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _5257_ (.A1(net335),
    .A2(net313),
    .B1(net263),
    .B2(net1650),
    .X(_0473_));
 sky130_fd_sc_hd__a22o_1 _5258_ (.A1(net337),
    .A2(net313),
    .B1(net263),
    .B2(net1084),
    .X(_0474_));
 sky130_fd_sc_hd__a22o_1 _5259_ (.A1(net357),
    .A2(net314),
    .B1(net264),
    .B2(net1572),
    .X(_0475_));
 sky130_fd_sc_hd__nor2_2 _5260_ (.A(_2654_),
    .B(_2661_),
    .Y(_2666_));
 sky130_fd_sc_hd__or2_1 _5261_ (.A(_2654_),
    .B(_2661_),
    .X(_2667_));
 sky130_fd_sc_hd__nor2_2 _5262_ (.A(net461),
    .B(net312),
    .Y(_2668_));
 sky130_fd_sc_hd__nand2_1 _5263_ (.A(net449),
    .B(_2667_),
    .Y(_2669_));
 sky130_fd_sc_hd__a22o_1 _5264_ (.A1(net356),
    .A2(net312),
    .B1(net262),
    .B2(net957),
    .X(_0476_));
 sky130_fd_sc_hd__o22a_1 _5265_ (.A1(_1689_),
    .A2(_2667_),
    .B1(_2669_),
    .B2(net905),
    .X(_0477_));
 sky130_fd_sc_hd__a22o_1 _5266_ (.A1(net329),
    .A2(net312),
    .B1(net262),
    .B2(net1666),
    .X(_0478_));
 sky130_fd_sc_hd__o22a_1 _5267_ (.A1(net330),
    .A2(_2667_),
    .B1(_2669_),
    .B2(net835),
    .X(_0479_));
 sky130_fd_sc_hd__a22o_1 _5268_ (.A1(net327),
    .A2(net311),
    .B1(net261),
    .B2(net1654),
    .X(_0480_));
 sky130_fd_sc_hd__a22o_1 _5269_ (.A1(net325),
    .A2(net312),
    .B1(net262),
    .B2(net1146),
    .X(_0481_));
 sky130_fd_sc_hd__a22o_1 _5270_ (.A1(net328),
    .A2(net312),
    .B1(net262),
    .B2(net1392),
    .X(_0482_));
 sky130_fd_sc_hd__a22o_1 _5271_ (.A1(net326),
    .A2(net311),
    .B1(net261),
    .B2(net1698),
    .X(_0483_));
 sky130_fd_sc_hd__a22o_1 _5272_ (.A1(net323),
    .A2(net312),
    .B1(net262),
    .B2(net1386),
    .X(_0484_));
 sky130_fd_sc_hd__a22o_1 _5273_ (.A1(net321),
    .A2(net312),
    .B1(net262),
    .B2(net1570),
    .X(_0485_));
 sky130_fd_sc_hd__a22o_1 _5274_ (.A1(net324),
    .A2(net312),
    .B1(net262),
    .B2(net1202),
    .X(_0486_));
 sky130_fd_sc_hd__a22o_1 _5275_ (.A1(net322),
    .A2(net311),
    .B1(net261),
    .B2(net1428),
    .X(_0487_));
 sky130_fd_sc_hd__a22o_1 _5276_ (.A1(net319),
    .A2(net312),
    .B1(net262),
    .B2(net1270),
    .X(_0488_));
 sky130_fd_sc_hd__a22o_1 _5277_ (.A1(net317),
    .A2(net312),
    .B1(net262),
    .B2(net1584),
    .X(_0489_));
 sky130_fd_sc_hd__a22o_1 _5278_ (.A1(net320),
    .A2(net312),
    .B1(net262),
    .B2(net1528),
    .X(_0490_));
 sky130_fd_sc_hd__a22o_1 _5279_ (.A1(net318),
    .A2(net311),
    .B1(net261),
    .B2(net1234),
    .X(_0491_));
 sky130_fd_sc_hd__a22o_1 _5280_ (.A1(net341),
    .A2(net311),
    .B1(net261),
    .B2(net1128),
    .X(_0492_));
 sky130_fd_sc_hd__a22o_1 _5281_ (.A1(net340),
    .A2(net312),
    .B1(net262),
    .B2(net1642),
    .X(_0493_));
 sky130_fd_sc_hd__a22o_1 _5282_ (.A1(net339),
    .A2(net311),
    .B1(net261),
    .B2(net1182),
    .X(_0494_));
 sky130_fd_sc_hd__a22o_1 _5283_ (.A1(net338),
    .A2(net311),
    .B1(net261),
    .B2(net1246),
    .X(_0495_));
 sky130_fd_sc_hd__a22o_1 _5284_ (.A1(net333),
    .A2(net311),
    .B1(net261),
    .B2(net1126),
    .X(_0496_));
 sky130_fd_sc_hd__a22o_1 _5285_ (.A1(net331),
    .A2(net312),
    .B1(net262),
    .B2(net1416),
    .X(_0497_));
 sky130_fd_sc_hd__a22o_1 _5286_ (.A1(net334),
    .A2(net311),
    .B1(net261),
    .B2(net1396),
    .X(_0498_));
 sky130_fd_sc_hd__a22o_1 _5287_ (.A1(net332),
    .A2(net311),
    .B1(net261),
    .B2(net1420),
    .X(_0499_));
 sky130_fd_sc_hd__a22o_1 _5288_ (.A1(net343),
    .A2(net311),
    .B1(net261),
    .B2(net1284),
    .X(_0500_));
 sky130_fd_sc_hd__a22o_1 _5289_ (.A1(net348),
    .A2(net312),
    .B1(net262),
    .B2(net977),
    .X(_0501_));
 sky130_fd_sc_hd__a22o_1 _5290_ (.A1(net344),
    .A2(net311),
    .B1(net261),
    .B2(net1168),
    .X(_0502_));
 sky130_fd_sc_hd__a22o_1 _5291_ (.A1(net342),
    .A2(net311),
    .B1(net261),
    .B2(net1350),
    .X(_0503_));
 sky130_fd_sc_hd__a22o_1 _5292_ (.A1(net336),
    .A2(net311),
    .B1(net261),
    .B2(net1352),
    .X(_0504_));
 sky130_fd_sc_hd__a22o_1 _5293_ (.A1(net335),
    .A2(net311),
    .B1(net261),
    .B2(net1662),
    .X(_0505_));
 sky130_fd_sc_hd__a22o_1 _5294_ (.A1(net337),
    .A2(net311),
    .B1(net261),
    .B2(net1124),
    .X(_0506_));
 sky130_fd_sc_hd__a22o_1 _5295_ (.A1(net357),
    .A2(net312),
    .B1(net262),
    .B2(net1466),
    .X(_0507_));
 sky130_fd_sc_hd__or3b_4 _5296_ (.A(_1407_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .C_N(_2653_),
    .X(_2670_));
 sky130_fd_sc_hd__nor2_2 _5297_ (.A(_2655_),
    .B(_2670_),
    .Y(_2671_));
 sky130_fd_sc_hd__or2_1 _5298_ (.A(_2655_),
    .B(_2670_),
    .X(_2672_));
 sky130_fd_sc_hd__nor2_2 _5299_ (.A(net466),
    .B(net309),
    .Y(_2673_));
 sky130_fd_sc_hd__nand2_1 _5300_ (.A(net450),
    .B(_2672_),
    .Y(_2674_));
 sky130_fd_sc_hd__o22a_1 _5301_ (.A1(net356),
    .A2(_2672_),
    .B1(_2674_),
    .B2(net869),
    .X(_0508_));
 sky130_fd_sc_hd__a22o_1 _5302_ (.A1(_1689_),
    .A2(net310),
    .B1(net260),
    .B2(net1068),
    .X(_0509_));
 sky130_fd_sc_hd__o22a_1 _5303_ (.A1(net329),
    .A2(_2672_),
    .B1(_2674_),
    .B2(net843),
    .X(_0510_));
 sky130_fd_sc_hd__o22a_1 _5304_ (.A1(net330),
    .A2(_2672_),
    .B1(_2674_),
    .B2(net965),
    .X(_0511_));
 sky130_fd_sc_hd__a22o_1 _5305_ (.A1(net327),
    .A2(net309),
    .B1(net259),
    .B2(net1330),
    .X(_0512_));
 sky130_fd_sc_hd__a22o_1 _5306_ (.A1(net325),
    .A2(net310),
    .B1(net260),
    .B2(net1388),
    .X(_0513_));
 sky130_fd_sc_hd__a22o_1 _5307_ (.A1(net328),
    .A2(net310),
    .B1(net260),
    .B2(net1470),
    .X(_0514_));
 sky130_fd_sc_hd__a22o_1 _5308_ (.A1(net326),
    .A2(net309),
    .B1(net259),
    .B2(net1772),
    .X(_0515_));
 sky130_fd_sc_hd__a22o_1 _5309_ (.A1(net323),
    .A2(net310),
    .B1(net260),
    .B2(net1026),
    .X(_0516_));
 sky130_fd_sc_hd__a22o_1 _5310_ (.A1(net321),
    .A2(net310),
    .B1(net260),
    .B2(net1634),
    .X(_0517_));
 sky130_fd_sc_hd__a22o_1 _5311_ (.A1(net324),
    .A2(net310),
    .B1(net260),
    .B2(net1018),
    .X(_0518_));
 sky130_fd_sc_hd__a22o_1 _5312_ (.A1(net322),
    .A2(net309),
    .B1(net259),
    .B2(net1003),
    .X(_0519_));
 sky130_fd_sc_hd__a22o_1 _5313_ (.A1(net319),
    .A2(net310),
    .B1(net260),
    .B2(net1682),
    .X(_0520_));
 sky130_fd_sc_hd__a22o_1 _5314_ (.A1(net317),
    .A2(net310),
    .B1(net260),
    .B2(net1520),
    .X(_0521_));
 sky130_fd_sc_hd__a22o_1 _5315_ (.A1(net320),
    .A2(net310),
    .B1(net260),
    .B2(net1512),
    .X(_0522_));
 sky130_fd_sc_hd__a22o_1 _5316_ (.A1(net318),
    .A2(net309),
    .B1(net259),
    .B2(net1116),
    .X(_0523_));
 sky130_fd_sc_hd__a22o_1 _5317_ (.A1(net341),
    .A2(net310),
    .B1(net259),
    .B2(net1198),
    .X(_0524_));
 sky130_fd_sc_hd__a22o_1 _5318_ (.A1(net340),
    .A2(net310),
    .B1(net260),
    .B2(net1600),
    .X(_0525_));
 sky130_fd_sc_hd__a22o_1 _5319_ (.A1(net339),
    .A2(net309),
    .B1(net259),
    .B2(net1232),
    .X(_0526_));
 sky130_fd_sc_hd__a22o_1 _5320_ (.A1(net338),
    .A2(net309),
    .B1(net259),
    .B2(net1562),
    .X(_0527_));
 sky130_fd_sc_hd__a22o_1 _5321_ (.A1(net333),
    .A2(net309),
    .B1(net259),
    .B2(net1690),
    .X(_0528_));
 sky130_fd_sc_hd__a22o_1 _5322_ (.A1(net331),
    .A2(net310),
    .B1(net260),
    .B2(net1076),
    .X(_0529_));
 sky130_fd_sc_hd__a22o_1 _5323_ (.A1(net334),
    .A2(net309),
    .B1(net259),
    .B2(net1298),
    .X(_0530_));
 sky130_fd_sc_hd__a22o_1 _5324_ (.A1(net332),
    .A2(net309),
    .B1(net259),
    .B2(net1506),
    .X(_0531_));
 sky130_fd_sc_hd__a22o_1 _5325_ (.A1(net343),
    .A2(net309),
    .B1(net259),
    .B2(net1318),
    .X(_0532_));
 sky130_fd_sc_hd__a22o_1 _5326_ (.A1(net348),
    .A2(net310),
    .B1(net260),
    .B2(net1382),
    .X(_0533_));
 sky130_fd_sc_hd__a22o_1 _5327_ (.A1(net344),
    .A2(net309),
    .B1(net259),
    .B2(net1554),
    .X(_0534_));
 sky130_fd_sc_hd__a22o_1 _5328_ (.A1(net342),
    .A2(net309),
    .B1(net259),
    .B2(net1502),
    .X(_0535_));
 sky130_fd_sc_hd__a22o_1 _5329_ (.A1(_1566_),
    .A2(net309),
    .B1(net259),
    .B2(net1590),
    .X(_0536_));
 sky130_fd_sc_hd__a22o_1 _5330_ (.A1(net335),
    .A2(net309),
    .B1(net259),
    .B2(net1015),
    .X(_0537_));
 sky130_fd_sc_hd__a22o_1 _5331_ (.A1(net337),
    .A2(net309),
    .B1(net259),
    .B2(net1136),
    .X(_0538_));
 sky130_fd_sc_hd__a22o_1 _5332_ (.A1(net357),
    .A2(net310),
    .B1(net260),
    .B2(net1092),
    .X(_0539_));
 sky130_fd_sc_hd__nor2_2 _5333_ (.A(_2655_),
    .B(_2660_),
    .Y(_2675_));
 sky130_fd_sc_hd__or2_2 _5334_ (.A(_2655_),
    .B(_2660_),
    .X(_2676_));
 sky130_fd_sc_hd__nor2_2 _5335_ (.A(net466),
    .B(net308),
    .Y(_2677_));
 sky130_fd_sc_hd__nand2_2 _5336_ (.A(net450),
    .B(_2676_),
    .Y(_2678_));
 sky130_fd_sc_hd__o22a_1 _5337_ (.A1(net356),
    .A2(_2676_),
    .B1(_2678_),
    .B2(net833),
    .X(_0540_));
 sky130_fd_sc_hd__o22a_1 _5338_ (.A1(_1689_),
    .A2(_2676_),
    .B1(_2678_),
    .B2(net851),
    .X(_0541_));
 sky130_fd_sc_hd__o22a_1 _5339_ (.A1(net329),
    .A2(_2676_),
    .B1(_2678_),
    .B2(net863),
    .X(_0542_));
 sky130_fd_sc_hd__o22a_1 _5340_ (.A1(net330),
    .A2(_2676_),
    .B1(_2678_),
    .B2(net895),
    .X(_0543_));
 sky130_fd_sc_hd__a22o_1 _5341_ (.A1(net327),
    .A2(net307),
    .B1(net257),
    .B2(net1660),
    .X(_0544_));
 sky130_fd_sc_hd__a22o_1 _5342_ (.A1(net325),
    .A2(net308),
    .B1(net258),
    .B2(net1524),
    .X(_0545_));
 sky130_fd_sc_hd__a22o_1 _5343_ (.A1(net328),
    .A2(net308),
    .B1(net258),
    .B2(net1228),
    .X(_0546_));
 sky130_fd_sc_hd__a22o_1 _5344_ (.A1(net326),
    .A2(net307),
    .B1(net257),
    .B2(net1564),
    .X(_0547_));
 sky130_fd_sc_hd__a22o_1 _5345_ (.A1(net323),
    .A2(net308),
    .B1(net258),
    .B2(net1644),
    .X(_0548_));
 sky130_fd_sc_hd__a22o_1 _5346_ (.A1(net321),
    .A2(net308),
    .B1(net258),
    .B2(net1020),
    .X(_0549_));
 sky130_fd_sc_hd__a22o_1 _5347_ (.A1(net324),
    .A2(net308),
    .B1(net258),
    .B2(net1504),
    .X(_0550_));
 sky130_fd_sc_hd__a22o_1 _5348_ (.A1(net322),
    .A2(net307),
    .B1(net257),
    .B2(net1162),
    .X(_0551_));
 sky130_fd_sc_hd__a22o_1 _5349_ (.A1(net319),
    .A2(net308),
    .B1(net258),
    .B2(net1630),
    .X(_0552_));
 sky130_fd_sc_hd__a22o_1 _5350_ (.A1(net317),
    .A2(net308),
    .B1(net258),
    .B2(net1582),
    .X(_0553_));
 sky130_fd_sc_hd__a22o_1 _5351_ (.A1(net320),
    .A2(net308),
    .B1(net258),
    .B2(net1480),
    .X(_0554_));
 sky130_fd_sc_hd__a22o_1 _5352_ (.A1(net318),
    .A2(net307),
    .B1(net257),
    .B2(net1166),
    .X(_0555_));
 sky130_fd_sc_hd__a22o_1 _5353_ (.A1(net341),
    .A2(net307),
    .B1(net257),
    .B2(net1007),
    .X(_0556_));
 sky130_fd_sc_hd__a22o_1 _5354_ (.A1(net340),
    .A2(net308),
    .B1(net258),
    .B2(net1412),
    .X(_0557_));
 sky130_fd_sc_hd__a22o_1 _5355_ (.A1(net339),
    .A2(net307),
    .B1(net257),
    .B2(net1172),
    .X(_0558_));
 sky130_fd_sc_hd__a22o_1 _5356_ (.A1(net338),
    .A2(net307),
    .B1(net257),
    .B2(net1304),
    .X(_0559_));
 sky130_fd_sc_hd__a22o_1 _5357_ (.A1(net333),
    .A2(net307),
    .B1(net257),
    .B2(net1354),
    .X(_0560_));
 sky130_fd_sc_hd__a22o_1 _5358_ (.A1(net331),
    .A2(net308),
    .B1(net258),
    .B2(net1046),
    .X(_0561_));
 sky130_fd_sc_hd__a22o_1 _5359_ (.A1(net334),
    .A2(net307),
    .B1(net257),
    .B2(net1550),
    .X(_0562_));
 sky130_fd_sc_hd__a22o_1 _5360_ (.A1(net332),
    .A2(net307),
    .B1(net257),
    .B2(net1120),
    .X(_0563_));
 sky130_fd_sc_hd__a22o_1 _5361_ (.A1(net343),
    .A2(net307),
    .B1(net257),
    .B2(net1028),
    .X(_0564_));
 sky130_fd_sc_hd__a22o_1 _5362_ (.A1(net348),
    .A2(net308),
    .B1(net258),
    .B2(net1220),
    .X(_0565_));
 sky130_fd_sc_hd__a22o_1 _5363_ (.A1(net344),
    .A2(net307),
    .B1(net257),
    .B2(net1164),
    .X(_0566_));
 sky130_fd_sc_hd__a22o_1 _5364_ (.A1(net342),
    .A2(net307),
    .B1(net257),
    .B2(net1418),
    .X(_0567_));
 sky130_fd_sc_hd__a22o_1 _5365_ (.A1(net336),
    .A2(net307),
    .B1(net257),
    .B2(net1394),
    .X(_0568_));
 sky130_fd_sc_hd__a22o_1 _5366_ (.A1(net335),
    .A2(net307),
    .B1(net257),
    .B2(net1374),
    .X(_0569_));
 sky130_fd_sc_hd__a22o_1 _5367_ (.A1(net337),
    .A2(net307),
    .B1(net257),
    .B2(net1158),
    .X(_0570_));
 sky130_fd_sc_hd__a22o_1 _5368_ (.A1(net357),
    .A2(net308),
    .B1(net258),
    .B2(net1316),
    .X(_0571_));
 sky130_fd_sc_hd__and2_2 _5369_ (.A(net176),
    .B(net225),
    .X(_2679_));
 sky130_fd_sc_hd__nand2_1 _5370_ (.A(net172),
    .B(net221),
    .Y(_2680_));
 sky130_fd_sc_hd__or3_2 _5371_ (.A(net2145),
    .B(net1980),
    .C(net2127),
    .X(_2681_));
 sky130_fd_sc_hd__or2_1 _5372_ (.A(net2210),
    .B(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ),
    .X(_2682_));
 sky130_fd_sc_hd__nor2_1 _5373_ (.A(_2177_),
    .B(net2211),
    .Y(_2683_));
 sky130_fd_sc_hd__or3_1 _5374_ (.A(_2177_),
    .B(_2681_),
    .C(net2211),
    .X(_2684_));
 sky130_fd_sc_hd__and3_1 _5375_ (.A(net176),
    .B(net225),
    .C(_2684_),
    .X(_2685_));
 sky130_fd_sc_hd__nand2_1 _5376_ (.A(net2170),
    .B(net2258),
    .Y(_2686_));
 sky130_fd_sc_hd__nor2_1 _5377_ (.A(net2211),
    .B(_2686_),
    .Y(_2687_));
 sky130_fd_sc_hd__and2b_1 _5378_ (.A_N(net1988),
    .B(_2687_),
    .X(_2688_));
 sky130_fd_sc_hd__a21o_1 _5379_ (.A1(_2681_),
    .A2(_2688_),
    .B1(_2683_),
    .X(_2689_));
 sky130_fd_sc_hd__and2b_1 _5380_ (.A_N(net2145),
    .B(_2689_),
    .X(_2690_));
 sky130_fd_sc_hd__nand2_1 _5381_ (.A(net2127),
    .B(_2690_),
    .Y(_2691_));
 sky130_fd_sc_hd__or2_1 _5382_ (.A(_1403_),
    .B(_2691_),
    .X(_2692_));
 sky130_fd_sc_hd__nand2_2 _5383_ (.A(net2145),
    .B(_2689_),
    .Y(_2693_));
 sky130_fd_sc_hd__o31a_1 _5384_ (.A1(net1980),
    .A2(net2127),
    .A3(_2693_),
    .B1(_2692_),
    .X(_2694_));
 sky130_fd_sc_hd__xnor2_1 _5385_ (.A(net1980),
    .B(net2127),
    .Y(_2695_));
 sky130_fd_sc_hd__nand2b_1 _5386_ (.A_N(_2695_),
    .B(_2690_),
    .Y(_2696_));
 sky130_fd_sc_hd__nor3_1 _5387_ (.A(net1988),
    .B(_2174_),
    .C(_2686_),
    .Y(_2697_));
 sky130_fd_sc_hd__or3_2 _5388_ (.A(net1988),
    .B(_2174_),
    .C(_2686_),
    .X(_2698_));
 sky130_fd_sc_hd__or3b_1 _5389_ (.A(_2174_),
    .B(net1988),
    .C_N(net2258),
    .X(_2699_));
 sky130_fd_sc_hd__o21ai_4 _5390_ (.A1(_2174_),
    .A2(_2177_),
    .B1(_2698_),
    .Y(_2700_));
 sky130_fd_sc_hd__nor3b_4 _5391_ (.A(net2258),
    .B(net2211),
    .C_N(net2170),
    .Y(_2701_));
 sky130_fd_sc_hd__or3b_1 _5392_ (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .B(_2682_),
    .C_N(net2170),
    .X(_2702_));
 sky130_fd_sc_hd__and2_1 _5393_ (.A(net1988),
    .B(_2701_),
    .X(_2703_));
 sky130_fd_sc_hd__nand2_1 _5394_ (.A(net1988),
    .B(_2701_),
    .Y(_2704_));
 sky130_fd_sc_hd__or4b_1 _5395_ (.A(_2689_),
    .B(_2700_),
    .C(_2703_),
    .D_N(_2176_),
    .X(_2705_));
 sky130_fd_sc_hd__and2_1 _5396_ (.A(_2696_),
    .B(_2705_),
    .X(_2706_));
 sky130_fd_sc_hd__o21bai_1 _5397_ (.A1(net1980),
    .A2(net2127),
    .B1_N(_2693_),
    .Y(_2707_));
 sky130_fd_sc_hd__o21a_1 _5398_ (.A1(net2145),
    .A2(_1403_),
    .B1(_2703_),
    .X(_2708_));
 sky130_fd_sc_hd__inv_2 _5399_ (.A(_2708_),
    .Y(_2709_));
 sky130_fd_sc_hd__o2111a_1 _5400_ (.A1(_0068_),
    .A2(_2697_),
    .B1(_2709_),
    .C1(_2692_),
    .D1(_2693_),
    .X(_2710_));
 sky130_fd_sc_hd__and3_1 _5401_ (.A(_2685_),
    .B(_2706_),
    .C(_2710_),
    .X(_0572_));
 sky130_fd_sc_hd__or2_1 _5402_ (.A(net1988),
    .B(net2171),
    .X(_2711_));
 sky130_fd_sc_hd__nor2_2 _5403_ (.A(net160),
    .B(_2711_),
    .Y(_0573_));
 sky130_fd_sc_hd__and3_2 _5404_ (.A(net2210),
    .B(net2254),
    .C(_2175_),
    .X(_2712_));
 sky130_fd_sc_hd__inv_2 _5405_ (.A(_2712_),
    .Y(_2713_));
 sky130_fd_sc_hd__and4bb_1 _5406_ (.A_N(_2683_),
    .B_N(_2688_),
    .C(_2713_),
    .D(_2679_),
    .X(_0574_));
 sky130_fd_sc_hd__nand2_4 _5407_ (.A(net1989),
    .B(_2713_),
    .Y(_2714_));
 sky130_fd_sc_hd__or3_1 _5408_ (.A(net1988),
    .B(net2170),
    .C(net2211),
    .X(_2715_));
 sky130_fd_sc_hd__nand2_1 _5409_ (.A(_2176_),
    .B(_2715_),
    .Y(_2716_));
 sky130_fd_sc_hd__o31a_1 _5410_ (.A1(_2687_),
    .A2(_2714_),
    .A3(_2716_),
    .B1(_2679_),
    .X(_0575_));
 sky130_fd_sc_hd__and3_1 _5411_ (.A(net925),
    .B(net176),
    .C(net227),
    .X(_0576_));
 sky130_fd_sc_hd__and3_1 _5412_ (.A(net1013),
    .B(net176),
    .C(net226),
    .X(_0577_));
 sky130_fd_sc_hd__and3_1 _5413_ (.A(net839),
    .B(net172),
    .C(net221),
    .X(_0578_));
 sky130_fd_sc_hd__and3_1 _5414_ (.A(net935),
    .B(net173),
    .C(net221),
    .X(_0579_));
 sky130_fd_sc_hd__and3_1 _5415_ (.A(net919),
    .B(net179),
    .C(net227),
    .X(_0580_));
 sky130_fd_sc_hd__and3_1 _5416_ (.A(net883),
    .B(net176),
    .C(net225),
    .X(_0581_));
 sky130_fd_sc_hd__and3_1 _5417_ (.A(net897),
    .B(net179),
    .C(net227),
    .X(_0582_));
 sky130_fd_sc_hd__and3_1 _5418_ (.A(net969),
    .B(net178),
    .C(net227),
    .X(_0583_));
 sky130_fd_sc_hd__and3_1 _5419_ (.A(net877),
    .B(net178),
    .C(net230),
    .X(_0584_));
 sky130_fd_sc_hd__and3_1 _5420_ (.A(net849),
    .B(net179),
    .C(net228),
    .X(_0585_));
 sky130_fd_sc_hd__and3_1 _5421_ (.A(net931),
    .B(net178),
    .C(net231),
    .X(_0586_));
 sky130_fd_sc_hd__and3_1 _5422_ (.A(net943),
    .B(net178),
    .C(net230),
    .X(_0587_));
 sky130_fd_sc_hd__and3_1 _5423_ (.A(net973),
    .B(net178),
    .C(net230),
    .X(_0588_));
 sky130_fd_sc_hd__and3_1 _5424_ (.A(net1152),
    .B(net169),
    .C(net214),
    .X(_0589_));
 sky130_fd_sc_hd__and3_1 _5425_ (.A(net921),
    .B(net169),
    .C(net214),
    .X(_0590_));
 sky130_fd_sc_hd__and3_1 _5426_ (.A(net951),
    .B(net169),
    .C(net215),
    .X(_0591_));
 sky130_fd_sc_hd__and3_1 _5427_ (.A(net985),
    .B(net173),
    .C(net217),
    .X(_0592_));
 sky130_fd_sc_hd__and3_1 _5428_ (.A(net1322),
    .B(net170),
    .C(net219),
    .X(_0593_));
 sky130_fd_sc_hd__and3_1 _5429_ (.A(net809),
    .B(net171),
    .C(net218),
    .X(_0594_));
 sky130_fd_sc_hd__and3_1 _5430_ (.A(net783),
    .B(net170),
    .C(net216),
    .X(_0595_));
 sky130_fd_sc_hd__and3_1 _5431_ (.A(net803),
    .B(net169),
    .C(net214),
    .X(_0596_));
 sky130_fd_sc_hd__and3_1 _5432_ (.A(net821),
    .B(net169),
    .C(net215),
    .X(_0597_));
 sky130_fd_sc_hd__and3_1 _5433_ (.A(net901),
    .B(net171),
    .C(net218),
    .X(_0598_));
 sky130_fd_sc_hd__and3_1 _5434_ (.A(net703),
    .B(net171),
    .C(net217),
    .X(_0599_));
 sky130_fd_sc_hd__and3_1 _5435_ (.A(net893),
    .B(net171),
    .C(net217),
    .X(_0600_));
 sky130_fd_sc_hd__and3_1 _5436_ (.A(net945),
    .B(net172),
    .C(net220),
    .X(_0601_));
 sky130_fd_sc_hd__and3_1 _5437_ (.A(net913),
    .B(net172),
    .C(net221),
    .X(_0602_));
 sky130_fd_sc_hd__and3_1 _5438_ (.A(net955),
    .B(net172),
    .C(net222),
    .X(_0603_));
 sky130_fd_sc_hd__and3_1 _5439_ (.A(net989),
    .B(net172),
    .C(net222),
    .X(_0604_));
 sky130_fd_sc_hd__and3_1 _5440_ (.A(net941),
    .B(net173),
    .C(net221),
    .X(_0605_));
 sky130_fd_sc_hd__and3_1 _5441_ (.A(net887),
    .B(net176),
    .C(net225),
    .X(_0606_));
 sky130_fd_sc_hd__and3_1 _5442_ (.A(net873),
    .B(net176),
    .C(net226),
    .X(_0607_));
 sky130_fd_sc_hd__and3_1 _5443_ (.A(net819),
    .B(net173),
    .C(net221),
    .X(_0608_));
 sky130_fd_sc_hd__and3_1 _5444_ (.A(net827),
    .B(net176),
    .C(net225),
    .X(_0609_));
 sky130_fd_sc_hd__and3_1 _5445_ (.A(net1130),
    .B(net176),
    .C(net225),
    .X(_0610_));
 sky130_fd_sc_hd__and3_1 _5446_ (.A(net875),
    .B(net176),
    .C(net225),
    .X(_0611_));
 sky130_fd_sc_hd__and3_1 _5447_ (.A(net853),
    .B(net179),
    .C(net227),
    .X(_0612_));
 sky130_fd_sc_hd__and3_1 _5448_ (.A(net823),
    .B(net178),
    .C(net230),
    .X(_0613_));
 sky130_fd_sc_hd__and3_1 _5449_ (.A(net961),
    .B(net178),
    .C(net227),
    .X(_0614_));
 sky130_fd_sc_hd__and3_1 _5450_ (.A(net987),
    .B(net178),
    .C(net230),
    .X(_0615_));
 sky130_fd_sc_hd__and3_1 _5451_ (.A(net937),
    .B(net179),
    .C(net231),
    .X(_0616_));
 sky130_fd_sc_hd__and3_1 _5452_ (.A(net899),
    .B(net178),
    .C(net230),
    .X(_0617_));
 sky130_fd_sc_hd__and3_1 _5453_ (.A(net967),
    .B(net178),
    .C(net230),
    .X(_0618_));
 sky130_fd_sc_hd__and3_1 _5454_ (.A(net995),
    .B(net169),
    .C(net214),
    .X(_0619_));
 sky130_fd_sc_hd__and3_1 _5455_ (.A(net979),
    .B(net169),
    .C(net216),
    .X(_0620_));
 sky130_fd_sc_hd__and3_1 _5456_ (.A(net993),
    .B(net170),
    .C(net219),
    .X(_0621_));
 sky130_fd_sc_hd__and3_1 _5457_ (.A(net813),
    .B(net169),
    .C(net216),
    .X(_0622_));
 sky130_fd_sc_hd__and3_1 _5458_ (.A(net1104),
    .B(net171),
    .C(net217),
    .X(_0623_));
 sky130_fd_sc_hd__and3_1 _5459_ (.A(net915),
    .B(net169),
    .C(net215),
    .X(_0624_));
 sky130_fd_sc_hd__and3_1 _5460_ (.A(net648),
    .B(net171),
    .C(net217),
    .X(_0625_));
 sky130_fd_sc_hd__and3_1 _5461_ (.A(net855),
    .B(net170),
    .C(net216),
    .X(_0626_));
 sky130_fd_sc_hd__and3_1 _5462_ (.A(net929),
    .B(net169),
    .C(net215),
    .X(_0627_));
 sky130_fd_sc_hd__and3_1 _5463_ (.A(net911),
    .B(net171),
    .C(net217),
    .X(_0628_));
 sky130_fd_sc_hd__and3_1 _5464_ (.A(net907),
    .B(net171),
    .C(net218),
    .X(_0629_));
 sky130_fd_sc_hd__and3_1 _5465_ (.A(net670),
    .B(net171),
    .C(net218),
    .X(_0630_));
 sky130_fd_sc_hd__and3_1 _5466_ (.A(net668),
    .B(net172),
    .C(net220),
    .X(_0631_));
 sky130_fd_sc_hd__and3_1 _5467_ (.A(net672),
    .B(net172),
    .C(net220),
    .X(_0632_));
 sky130_fd_sc_hd__and3_1 _5468_ (.A(net1098),
    .B(net172),
    .C(net220),
    .X(_0633_));
 sky130_fd_sc_hd__and3_1 _5469_ (.A(net933),
    .B(net172),
    .C(net221),
    .X(_0634_));
 sky130_fd_sc_hd__and3_1 _5470_ (.A(net1310),
    .B(net172),
    .C(net222),
    .X(_0635_));
 sky130_fd_sc_hd__nor2_1 _5471_ (.A(_1402_),
    .B(net160),
    .Y(_0636_));
 sky130_fd_sc_hd__and3_1 _5472_ (.A(net385),
    .B(net177),
    .C(net228),
    .X(_0637_));
 sky130_fd_sc_hd__and3_1 _5473_ (.A(net375),
    .B(net177),
    .C(net229),
    .X(_0638_));
 sky130_fd_sc_hd__and3_1 _5474_ (.A(net369),
    .B(net177),
    .C(net228),
    .X(_0639_));
 sky130_fd_sc_hd__and3_1 _5475_ (.A(net424),
    .B(net177),
    .C(net229),
    .X(_0640_));
 sky130_fd_sc_hd__and3_1 _5476_ (.A(net414),
    .B(net177),
    .C(net229),
    .X(_0641_));
 sky130_fd_sc_hd__and3_1 _5477_ (.A(net404),
    .B(net177),
    .C(net229),
    .X(_0642_));
 sky130_fd_sc_hd__and3_1 _5478_ (.A(net399),
    .B(net179),
    .C(net229),
    .X(_0643_));
 sky130_fd_sc_hd__and3_1 _5479_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[0] ),
    .B(net177),
    .C(net228),
    .X(_0644_));
 sky130_fd_sc_hd__and3_1 _5480_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[1] ),
    .B(net177),
    .C(net228),
    .X(_0645_));
 sky130_fd_sc_hd__and3_1 _5481_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[2] ),
    .B(net174),
    .C(net223),
    .X(_0646_));
 sky130_fd_sc_hd__and3_1 _5482_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[3] ),
    .B(net174),
    .C(net223),
    .X(_0647_));
 sky130_fd_sc_hd__and3_1 _5483_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[4] ),
    .B(net170),
    .C(net216),
    .X(_0648_));
 sky130_fd_sc_hd__and3_1 _5484_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[5] ),
    .B(net174),
    .C(net223),
    .X(_0649_));
 sky130_fd_sc_hd__and3_1 _5485_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[6] ),
    .B(net175),
    .C(net224),
    .X(_0650_));
 sky130_fd_sc_hd__and3_1 _5486_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[7] ),
    .B(net168),
    .C(net212),
    .X(_0651_));
 sky130_fd_sc_hd__and3_1 _5487_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[8] ),
    .B(net177),
    .C(net228),
    .X(_0652_));
 sky130_fd_sc_hd__and3_1 _5488_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[9] ),
    .B(net175),
    .C(net224),
    .X(_0653_));
 sky130_fd_sc_hd__and3_1 _5489_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[10] ),
    .B(net175),
    .C(net224),
    .X(_0654_));
 sky130_fd_sc_hd__and3_1 _5490_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[11] ),
    .B(net168),
    .C(net212),
    .X(_0655_));
 sky130_fd_sc_hd__and3_1 _5491_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[12] ),
    .B(net175),
    .C(net224),
    .X(_0656_));
 sky130_fd_sc_hd__and3_1 _5492_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[13] ),
    .B(net174),
    .C(net223),
    .X(_0657_));
 sky130_fd_sc_hd__and3_1 _5493_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[14] ),
    .B(net174),
    .C(net223),
    .X(_0658_));
 sky130_fd_sc_hd__and3_1 _5494_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[15] ),
    .B(net167),
    .C(net213),
    .X(_0659_));
 sky130_fd_sc_hd__and3_1 _5495_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[16] ),
    .B(net167),
    .C(net212),
    .X(_0660_));
 sky130_fd_sc_hd__and3_1 _5496_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[17] ),
    .B(net174),
    .C(net228),
    .X(_0661_));
 sky130_fd_sc_hd__and3_1 _5497_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[18] ),
    .B(net167),
    .C(net213),
    .X(_0662_));
 sky130_fd_sc_hd__and3_1 _5498_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[19] ),
    .B(net168),
    .C(net212),
    .X(_0663_));
 sky130_fd_sc_hd__and3_1 _5499_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[20] ),
    .B(net167),
    .C(net213),
    .X(_0664_));
 sky130_fd_sc_hd__and3_1 _5500_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[21] ),
    .B(net174),
    .C(net223),
    .X(_0665_));
 sky130_fd_sc_hd__and3_1 _5501_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[22] ),
    .B(net168),
    .C(net213),
    .X(_0666_));
 sky130_fd_sc_hd__and3_1 _5502_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[23] ),
    .B(net167),
    .C(net213),
    .X(_0667_));
 sky130_fd_sc_hd__and3_1 _5503_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[24] ),
    .B(net169),
    .C(net216),
    .X(_0668_));
 sky130_fd_sc_hd__and3_1 _5504_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[25] ),
    .B(net167),
    .C(net212),
    .X(_0669_));
 sky130_fd_sc_hd__and3_1 _5505_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[26] ),
    .B(net167),
    .C(net213),
    .X(_0670_));
 sky130_fd_sc_hd__and3_1 _5506_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[27] ),
    .B(net167),
    .C(net213),
    .X(_0671_));
 sky130_fd_sc_hd__and3_1 _5507_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[28] ),
    .B(net168),
    .C(net212),
    .X(_0672_));
 sky130_fd_sc_hd__and3_1 _5508_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[29] ),
    .B(net170),
    .C(net216),
    .X(_0673_));
 sky130_fd_sc_hd__and3_1 _5509_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[30] ),
    .B(net168),
    .C(net212),
    .X(_0674_));
 sky130_fd_sc_hd__and3_1 _5510_ (.A(\U_DATAPATH.U_ID_EX.i_rs2_ID[31] ),
    .B(net174),
    .C(net212),
    .X(_0675_));
 sky130_fd_sc_hd__and3_1 _5511_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[0] ),
    .B(net179),
    .C(net228),
    .X(_0676_));
 sky130_fd_sc_hd__and3_1 _5512_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[1] ),
    .B(net174),
    .C(net224),
    .X(_0677_));
 sky130_fd_sc_hd__and3_1 _5513_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[2] ),
    .B(net174),
    .C(net223),
    .X(_0678_));
 sky130_fd_sc_hd__and3_1 _5514_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[3] ),
    .B(net175),
    .C(net223),
    .X(_0679_));
 sky130_fd_sc_hd__and3_1 _5515_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[4] ),
    .B(net167),
    .C(net216),
    .X(_0680_));
 sky130_fd_sc_hd__and3_1 _5516_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[5] ),
    .B(net174),
    .C(net223),
    .X(_0681_));
 sky130_fd_sc_hd__and3_1 _5517_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[6] ),
    .B(net175),
    .C(net224),
    .X(_0682_));
 sky130_fd_sc_hd__and3_1 _5518_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[7] ),
    .B(net168),
    .C(net232),
    .X(_0683_));
 sky130_fd_sc_hd__and3_1 _5519_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[8] ),
    .B(net177),
    .C(net228),
    .X(_0684_));
 sky130_fd_sc_hd__and3_1 _5520_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[9] ),
    .B(net175),
    .C(net224),
    .X(_0685_));
 sky130_fd_sc_hd__and3_1 _5521_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[10] ),
    .B(net175),
    .C(net224),
    .X(_0686_));
 sky130_fd_sc_hd__and3_1 _5522_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[11] ),
    .B(net168),
    .C(net212),
    .X(_0687_));
 sky130_fd_sc_hd__and3_1 _5523_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[12] ),
    .B(net175),
    .C(net224),
    .X(_0688_));
 sky130_fd_sc_hd__and3_1 _5524_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[13] ),
    .B(net174),
    .C(net223),
    .X(_0689_));
 sky130_fd_sc_hd__and3_1 _5525_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[14] ),
    .B(net174),
    .C(net223),
    .X(_0690_));
 sky130_fd_sc_hd__and3_1 _5526_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[15] ),
    .B(net167),
    .C(net212),
    .X(_0691_));
 sky130_fd_sc_hd__and3_1 _5527_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[16] ),
    .B(net174),
    .C(net212),
    .X(_0692_));
 sky130_fd_sc_hd__and3_1 _5528_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[17] ),
    .B(net175),
    .C(net223),
    .X(_0693_));
 sky130_fd_sc_hd__and3_1 _5529_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[18] ),
    .B(net167),
    .C(net213),
    .X(_0694_));
 sky130_fd_sc_hd__and3_1 _5530_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[19] ),
    .B(net168),
    .C(net212),
    .X(_0695_));
 sky130_fd_sc_hd__and3_1 _5531_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[20] ),
    .B(net167),
    .C(net213),
    .X(_0696_));
 sky130_fd_sc_hd__and3_1 _5532_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[21] ),
    .B(net174),
    .C(net223),
    .X(_0697_));
 sky130_fd_sc_hd__and3_1 _5533_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[22] ),
    .B(net168),
    .C(net212),
    .X(_0698_));
 sky130_fd_sc_hd__and3_1 _5534_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[23] ),
    .B(net167),
    .C(net213),
    .X(_0699_));
 sky130_fd_sc_hd__and3_1 _5535_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[24] ),
    .B(net170),
    .C(net216),
    .X(_0700_));
 sky130_fd_sc_hd__and3_1 _5536_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[25] ),
    .B(net167),
    .C(net212),
    .X(_0701_));
 sky130_fd_sc_hd__and3_1 _5537_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[26] ),
    .B(net167),
    .C(net213),
    .X(_0702_));
 sky130_fd_sc_hd__and3_1 _5538_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[27] ),
    .B(net167),
    .C(net213),
    .X(_0703_));
 sky130_fd_sc_hd__and3_1 _5539_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[28] ),
    .B(net168),
    .C(net212),
    .X(_0704_));
 sky130_fd_sc_hd__and3_1 _5540_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[29] ),
    .B(net170),
    .C(net216),
    .X(_0705_));
 sky130_fd_sc_hd__and3_1 _5541_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[30] ),
    .B(net168),
    .C(net212),
    .X(_0706_));
 sky130_fd_sc_hd__and3_1 _5542_ (.A(\U_DATAPATH.U_ID_EX.i_rs1_ID[31] ),
    .B(net174),
    .C(net223),
    .X(_0707_));
 sky130_fd_sc_hd__nor2_1 _5543_ (.A(net1958),
    .B(net160),
    .Y(_0708_));
 sky130_fd_sc_hd__and3_1 _5544_ (.A(net1991),
    .B(net177),
    .C(net229),
    .X(_0709_));
 sky130_fd_sc_hd__and3_1 _5545_ (.A(net2121),
    .B(net177),
    .C(net228),
    .X(_0710_));
 sky130_fd_sc_hd__and3_1 _5546_ (.A(net2118),
    .B(net177),
    .C(net229),
    .X(_0711_));
 sky130_fd_sc_hd__nor2_1 _5547_ (.A(net160),
    .B(_2704_),
    .Y(_0712_));
 sky130_fd_sc_hd__nor2_1 _5548_ (.A(net160),
    .B(_2713_),
    .Y(_0713_));
 sky130_fd_sc_hd__and2_1 _5549_ (.A(net458),
    .B(net953),
    .X(_0714_));
 sky130_fd_sc_hd__and2_1 _5550_ (.A(net453),
    .B(net927),
    .X(_0715_));
 sky130_fd_sc_hd__and2_1 _5551_ (.A(net451),
    .B(_1913_),
    .X(_0716_));
 sky130_fd_sc_hd__and2_1 _5552_ (.A(net452),
    .B(net2132),
    .X(_0717_));
 sky130_fd_sc_hd__and2_1 _5553_ (.A(net441),
    .B(net2205),
    .X(_0718_));
 sky130_fd_sc_hd__and2_1 _5554_ (.A(net452),
    .B(net2209),
    .X(_0719_));
 sky130_fd_sc_hd__and2_1 _5555_ (.A(net452),
    .B(net2245),
    .X(_0720_));
 sky130_fd_sc_hd__and2_1 _5556_ (.A(net452),
    .B(net2219),
    .X(_0721_));
 sky130_fd_sc_hd__and2_1 _5557_ (.A(net451),
    .B(net2143),
    .X(_0722_));
 sky130_fd_sc_hd__and2_1 _5558_ (.A(net451),
    .B(net2234),
    .X(_0723_));
 sky130_fd_sc_hd__and2_1 _5559_ (.A(net455),
    .B(net2287),
    .X(_0724_));
 sky130_fd_sc_hd__and2_1 _5560_ (.A(net453),
    .B(net2055),
    .X(_0725_));
 sky130_fd_sc_hd__and2_1 _5561_ (.A(net455),
    .B(net2333),
    .X(_0726_));
 sky130_fd_sc_hd__and2_1 _5562_ (.A(net456),
    .B(net2187),
    .X(_0727_));
 sky130_fd_sc_hd__and2_1 _5563_ (.A(net455),
    .B(net2166),
    .X(_0728_));
 sky130_fd_sc_hd__and2_1 _5564_ (.A(net436),
    .B(net2063),
    .X(_0729_));
 sky130_fd_sc_hd__and2_1 _5565_ (.A(net435),
    .B(net2215),
    .X(_0730_));
 sky130_fd_sc_hd__and2_1 _5566_ (.A(net436),
    .B(net2043),
    .X(_0731_));
 sky130_fd_sc_hd__and2_1 _5567_ (.A(net440),
    .B(net2015),
    .X(_0732_));
 sky130_fd_sc_hd__and2_1 _5568_ (.A(net437),
    .B(net2180),
    .X(_0733_));
 sky130_fd_sc_hd__and2_1 _5569_ (.A(net438),
    .B(net2326),
    .X(_0734_));
 sky130_fd_sc_hd__and2_1 _5570_ (.A(net443),
    .B(net2279),
    .X(_0735_));
 sky130_fd_sc_hd__and2_1 _5571_ (.A(net437),
    .B(net2230),
    .X(_0736_));
 sky130_fd_sc_hd__nor2_1 _5572_ (.A(net463),
    .B(net2273),
    .Y(_0737_));
 sky130_fd_sc_hd__and2_1 _5573_ (.A(net439),
    .B(net2154),
    .X(_0738_));
 sky130_fd_sc_hd__nor2_1 _5574_ (.A(net463),
    .B(net2312),
    .Y(_0739_));
 sky130_fd_sc_hd__and2_1 _5575_ (.A(net439),
    .B(net2226),
    .X(_0740_));
 sky130_fd_sc_hd__and2_1 _5576_ (.A(net440),
    .B(net2197),
    .X(_0741_));
 sky130_fd_sc_hd__and2_1 _5577_ (.A(net441),
    .B(net2202),
    .X(_0742_));
 sky130_fd_sc_hd__and2_1 _5578_ (.A(net442),
    .B(net2032),
    .X(_0743_));
 sky130_fd_sc_hd__and2_1 _5579_ (.A(net441),
    .B(net2252),
    .X(_0744_));
 sky130_fd_sc_hd__and2_1 _5580_ (.A(net441),
    .B(net2027),
    .X(_0745_));
 sky130_fd_sc_hd__or2_4 _5581_ (.A(_1409_),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .X(_2717_));
 sky130_fd_sc_hd__nor2_2 _5582_ (.A(_2660_),
    .B(_2717_),
    .Y(_2718_));
 sky130_fd_sc_hd__or2_2 _5583_ (.A(_2660_),
    .B(_2717_),
    .X(_2719_));
 sky130_fd_sc_hd__nor2_2 _5584_ (.A(net466),
    .B(net306),
    .Y(_2720_));
 sky130_fd_sc_hd__nand2_1 _5585_ (.A(net449),
    .B(_2719_),
    .Y(_2721_));
 sky130_fd_sc_hd__o22a_1 _5586_ (.A1(net356),
    .A2(_2719_),
    .B1(_2721_),
    .B2(net917),
    .X(_0746_));
 sky130_fd_sc_hd__o22a_1 _5587_ (.A1(_1689_),
    .A2(_2719_),
    .B1(_2721_),
    .B2(net845),
    .X(_0747_));
 sky130_fd_sc_hd__o22a_1 _5588_ (.A1(net329),
    .A2(_2719_),
    .B1(_2721_),
    .B2(net865),
    .X(_0748_));
 sky130_fd_sc_hd__a22o_1 _5589_ (.A1(net330),
    .A2(net306),
    .B1(net256),
    .B2(net1604),
    .X(_0749_));
 sky130_fd_sc_hd__a22o_1 _5590_ (.A1(net327),
    .A2(net305),
    .B1(net255),
    .B2(net1332),
    .X(_0750_));
 sky130_fd_sc_hd__a22o_1 _5591_ (.A1(net325),
    .A2(net306),
    .B1(net256),
    .B2(net1108),
    .X(_0751_));
 sky130_fd_sc_hd__a22o_1 _5592_ (.A1(net328),
    .A2(net306),
    .B1(net256),
    .B2(net997),
    .X(_0752_));
 sky130_fd_sc_hd__a22o_1 _5593_ (.A1(net326),
    .A2(net305),
    .B1(net255),
    .B2(net1534),
    .X(_0753_));
 sky130_fd_sc_hd__a22o_1 _5594_ (.A1(net323),
    .A2(net306),
    .B1(net256),
    .B2(net1256),
    .X(_0754_));
 sky130_fd_sc_hd__a22o_1 _5595_ (.A1(net321),
    .A2(net306),
    .B1(net256),
    .B2(net1118),
    .X(_0755_));
 sky130_fd_sc_hd__a22o_1 _5596_ (.A1(net324),
    .A2(net306),
    .B1(net256),
    .B2(net1390),
    .X(_0756_));
 sky130_fd_sc_hd__a22o_1 _5597_ (.A1(net322),
    .A2(net305),
    .B1(net255),
    .B2(net1370),
    .X(_0757_));
 sky130_fd_sc_hd__a22o_1 _5598_ (.A1(net319),
    .A2(net306),
    .B1(net256),
    .B2(net1216),
    .X(_0758_));
 sky130_fd_sc_hd__a22o_1 _5599_ (.A1(net317),
    .A2(net306),
    .B1(net256),
    .B2(net1758),
    .X(_0759_));
 sky130_fd_sc_hd__a22o_1 _5600_ (.A1(net320),
    .A2(net306),
    .B1(net256),
    .B2(net1260),
    .X(_0760_));
 sky130_fd_sc_hd__a22o_1 _5601_ (.A1(net318),
    .A2(net305),
    .B1(net255),
    .B2(net1062),
    .X(_0761_));
 sky130_fd_sc_hd__a22o_1 _5602_ (.A1(net341),
    .A2(net306),
    .B1(net256),
    .B2(net1384),
    .X(_0762_));
 sky130_fd_sc_hd__a22o_1 _5603_ (.A1(net340),
    .A2(net306),
    .B1(net256),
    .B2(net1490),
    .X(_0763_));
 sky130_fd_sc_hd__a22o_1 _5604_ (.A1(net339),
    .A2(net305),
    .B1(net255),
    .B2(net1100),
    .X(_0764_));
 sky130_fd_sc_hd__a22o_1 _5605_ (.A1(net338),
    .A2(net305),
    .B1(net255),
    .B2(net1344),
    .X(_0765_));
 sky130_fd_sc_hd__a22o_1 _5606_ (.A1(net333),
    .A2(net305),
    .B1(net255),
    .B2(net1070),
    .X(_0766_));
 sky130_fd_sc_hd__a22o_1 _5607_ (.A1(net331),
    .A2(net306),
    .B1(net256),
    .B2(net1288),
    .X(_0767_));
 sky130_fd_sc_hd__a22o_1 _5608_ (.A1(net334),
    .A2(net305),
    .B1(net255),
    .B2(net1710),
    .X(_0768_));
 sky130_fd_sc_hd__a22o_1 _5609_ (.A1(net332),
    .A2(net305),
    .B1(net255),
    .B2(net1144),
    .X(_0769_));
 sky130_fd_sc_hd__a22o_1 _5610_ (.A1(net343),
    .A2(net305),
    .B1(net255),
    .B2(net1678),
    .X(_0770_));
 sky130_fd_sc_hd__a22o_1 _5611_ (.A1(net348),
    .A2(net305),
    .B1(net255),
    .B2(net1484),
    .X(_0771_));
 sky130_fd_sc_hd__a22o_1 _5612_ (.A1(net344),
    .A2(net305),
    .B1(net255),
    .B2(net1112),
    .X(_0772_));
 sky130_fd_sc_hd__a22o_1 _5613_ (.A1(net342),
    .A2(net305),
    .B1(net255),
    .B2(net1366),
    .X(_0773_));
 sky130_fd_sc_hd__a22o_1 _5614_ (.A1(net336),
    .A2(net305),
    .B1(net255),
    .B2(net1436),
    .X(_0774_));
 sky130_fd_sc_hd__a22o_1 _5615_ (.A1(net335),
    .A2(net305),
    .B1(net255),
    .B2(net1680),
    .X(_0775_));
 sky130_fd_sc_hd__a22o_1 _5616_ (.A1(net337),
    .A2(net305),
    .B1(net255),
    .B2(net1552),
    .X(_0776_));
 sky130_fd_sc_hd__a22o_1 _5617_ (.A1(net357),
    .A2(net306),
    .B1(net256),
    .B2(net1294),
    .X(_0777_));
 sky130_fd_sc_hd__nor2_2 _5618_ (.A(_2661_),
    .B(_2670_),
    .Y(_2722_));
 sky130_fd_sc_hd__or2_1 _5619_ (.A(_2661_),
    .B(_2670_),
    .X(_2723_));
 sky130_fd_sc_hd__nor2_2 _5620_ (.A(net466),
    .B(net304),
    .Y(_2724_));
 sky130_fd_sc_hd__nand2_1 _5621_ (.A(net450),
    .B(_2723_),
    .Y(_2725_));
 sky130_fd_sc_hd__o22a_1 _5622_ (.A1(net356),
    .A2(_2723_),
    .B1(_2725_),
    .B2(net829),
    .X(_0778_));
 sky130_fd_sc_hd__a22o_1 _5623_ (.A1(_1689_),
    .A2(net304),
    .B1(net254),
    .B2(net1048),
    .X(_0779_));
 sky130_fd_sc_hd__a22o_1 _5624_ (.A1(net329),
    .A2(net304),
    .B1(net254),
    .B2(net1300),
    .X(_0780_));
 sky130_fd_sc_hd__o22a_1 _5625_ (.A1(net330),
    .A2(_2723_),
    .B1(_2725_),
    .B2(net881),
    .X(_0781_));
 sky130_fd_sc_hd__a22o_1 _5626_ (.A1(net327),
    .A2(net303),
    .B1(net253),
    .B2(net1194),
    .X(_0782_));
 sky130_fd_sc_hd__a22o_1 _5627_ (.A1(net325),
    .A2(net304),
    .B1(net254),
    .B2(net1430),
    .X(_0783_));
 sky130_fd_sc_hd__a22o_1 _5628_ (.A1(net328),
    .A2(net304),
    .B1(net254),
    .B2(net1264),
    .X(_0784_));
 sky130_fd_sc_hd__a22o_1 _5629_ (.A1(net326),
    .A2(net303),
    .B1(net253),
    .B2(net1608),
    .X(_0785_));
 sky130_fd_sc_hd__a22o_1 _5630_ (.A1(net323),
    .A2(net304),
    .B1(net254),
    .B2(net1096),
    .X(_0786_));
 sky130_fd_sc_hd__a22o_1 _5631_ (.A1(net321),
    .A2(net304),
    .B1(net254),
    .B2(net1640),
    .X(_0787_));
 sky130_fd_sc_hd__a22o_1 _5632_ (.A1(net324),
    .A2(net304),
    .B1(net254),
    .B2(net1138),
    .X(_0788_));
 sky130_fd_sc_hd__a22o_1 _5633_ (.A1(net322),
    .A2(net303),
    .B1(net253),
    .B2(net1516),
    .X(_0789_));
 sky130_fd_sc_hd__a22o_1 _5634_ (.A1(net319),
    .A2(net304),
    .B1(net254),
    .B2(net1036),
    .X(_0790_));
 sky130_fd_sc_hd__a22o_1 _5635_ (.A1(net317),
    .A2(net304),
    .B1(net254),
    .B2(net1440),
    .X(_0791_));
 sky130_fd_sc_hd__a22o_1 _5636_ (.A1(net320),
    .A2(net304),
    .B1(net254),
    .B2(net1170),
    .X(_0792_));
 sky130_fd_sc_hd__a22o_1 _5637_ (.A1(net318),
    .A2(net303),
    .B1(net253),
    .B2(net1424),
    .X(_0793_));
 sky130_fd_sc_hd__a22o_1 _5638_ (.A1(net341),
    .A2(net303),
    .B1(net253),
    .B2(net1434),
    .X(_0794_));
 sky130_fd_sc_hd__a22o_1 _5639_ (.A1(net340),
    .A2(net304),
    .B1(net254),
    .B2(net1566),
    .X(_0795_));
 sky130_fd_sc_hd__a22o_1 _5640_ (.A1(net339),
    .A2(net303),
    .B1(net253),
    .B2(net1005),
    .X(_0796_));
 sky130_fd_sc_hd__a22o_1 _5641_ (.A1(net338),
    .A2(net303),
    .B1(net253),
    .B2(net1494),
    .X(_0797_));
 sky130_fd_sc_hd__a22o_1 _5642_ (.A1(net333),
    .A2(net303),
    .B1(net253),
    .B2(net1042),
    .X(_0798_));
 sky130_fd_sc_hd__a22o_1 _5643_ (.A1(net331),
    .A2(net304),
    .B1(net254),
    .B2(net1102),
    .X(_0799_));
 sky130_fd_sc_hd__a22o_1 _5644_ (.A1(net334),
    .A2(net303),
    .B1(net253),
    .B2(net1368),
    .X(_0800_));
 sky130_fd_sc_hd__a22o_1 _5645_ (.A1(net332),
    .A2(net303),
    .B1(net253),
    .B2(net1266),
    .X(_0801_));
 sky130_fd_sc_hd__a22o_1 _5646_ (.A1(net343),
    .A2(net303),
    .B1(net253),
    .B2(net1476),
    .X(_0802_));
 sky130_fd_sc_hd__a22o_1 _5647_ (.A1(net348),
    .A2(net304),
    .B1(net254),
    .B2(net1001),
    .X(_0803_));
 sky130_fd_sc_hd__a22o_1 _5648_ (.A1(net344),
    .A2(net303),
    .B1(net253),
    .B2(net959),
    .X(_0804_));
 sky130_fd_sc_hd__a22o_1 _5649_ (.A1(net342),
    .A2(net303),
    .B1(net253),
    .B2(net1492),
    .X(_0805_));
 sky130_fd_sc_hd__a22o_1 _5650_ (.A1(net336),
    .A2(net303),
    .B1(net253),
    .B2(net1218),
    .X(_0806_));
 sky130_fd_sc_hd__a22o_1 _5651_ (.A1(net335),
    .A2(net303),
    .B1(net253),
    .B2(net1210),
    .X(_0807_));
 sky130_fd_sc_hd__a22o_1 _5652_ (.A1(net337),
    .A2(net303),
    .B1(net253),
    .B2(net1314),
    .X(_0808_));
 sky130_fd_sc_hd__a22o_1 _5653_ (.A1(net357),
    .A2(net304),
    .B1(net254),
    .B2(net1276),
    .X(_0809_));
 sky130_fd_sc_hd__and2_1 _5654_ (.A(net458),
    .B(net2102),
    .X(_0810_));
 sky130_fd_sc_hd__and2_1 _5655_ (.A(net454),
    .B(net2087),
    .X(_0811_));
 sky130_fd_sc_hd__and2_1 _5656_ (.A(net454),
    .B(net2136),
    .X(_0812_));
 sky130_fd_sc_hd__and2_1 _5657_ (.A(net458),
    .B(net861),
    .X(_0813_));
 sky130_fd_sc_hd__and2_1 _5658_ (.A(net452),
    .B(net707),
    .X(_0814_));
 sky130_fd_sc_hd__and2_1 _5659_ (.A(net452),
    .B(net719),
    .X(_0815_));
 sky130_fd_sc_hd__and2_1 _5660_ (.A(net441),
    .B(net640),
    .X(_0816_));
 sky130_fd_sc_hd__and2_1 _5661_ (.A(net442),
    .B(net723),
    .X(_0817_));
 sky130_fd_sc_hd__and2_1 _5662_ (.A(net451),
    .B(net721),
    .X(_0818_));
 sky130_fd_sc_hd__and2_1 _5663_ (.A(net452),
    .B(net815),
    .X(_0819_));
 sky130_fd_sc_hd__and2_1 _5664_ (.A(net451),
    .B(net749),
    .X(_0820_));
 sky130_fd_sc_hd__and2_1 _5665_ (.A(net451),
    .B(net753),
    .X(_0821_));
 sky130_fd_sc_hd__and2_1 _5666_ (.A(net455),
    .B(net690),
    .X(_0822_));
 sky130_fd_sc_hd__and2_1 _5667_ (.A(net458),
    .B(net735),
    .X(_0823_));
 sky130_fd_sc_hd__and2_1 _5668_ (.A(net457),
    .B(net731),
    .X(_0824_));
 sky130_fd_sc_hd__and2_1 _5669_ (.A(net456),
    .B(net757),
    .X(_0825_));
 sky130_fd_sc_hd__and2_1 _5670_ (.A(net455),
    .B(net654),
    .X(_0826_));
 sky130_fd_sc_hd__and2_1 _5671_ (.A(net435),
    .B(net682),
    .X(_0827_));
 sky130_fd_sc_hd__and2_1 _5672_ (.A(net435),
    .B(net777),
    .X(_0828_));
 sky130_fd_sc_hd__and2_1 _5673_ (.A(net436),
    .B(net709),
    .X(_0829_));
 sky130_fd_sc_hd__and2_1 _5674_ (.A(net439),
    .B(net807),
    .X(_0830_));
 sky130_fd_sc_hd__and2_1 _5675_ (.A(net437),
    .B(net811),
    .X(_0831_));
 sky130_fd_sc_hd__and2_1 _5676_ (.A(net438),
    .B(net711),
    .X(_0832_));
 sky130_fd_sc_hd__and2_1 _5677_ (.A(net437),
    .B(net622),
    .X(_0833_));
 sky130_fd_sc_hd__and2_1 _5678_ (.A(net438),
    .B(net632),
    .X(_0834_));
 sky130_fd_sc_hd__and2_1 _5679_ (.A(net436),
    .B(net805),
    .X(_0835_));
 sky130_fd_sc_hd__and2_1 _5680_ (.A(net439),
    .B(net727),
    .X(_0836_));
 sky130_fd_sc_hd__and2_1 _5681_ (.A(net440),
    .B(net759),
    .X(_0837_));
 sky130_fd_sc_hd__and2_1 _5682_ (.A(net439),
    .B(net684),
    .X(_0838_));
 sky130_fd_sc_hd__and2_1 _5683_ (.A(net440),
    .B(net755),
    .X(_0839_));
 sky130_fd_sc_hd__and2_1 _5684_ (.A(net441),
    .B(net656),
    .X(_0840_));
 sky130_fd_sc_hd__and2_1 _5685_ (.A(net440),
    .B(net747),
    .X(_0841_));
 sky130_fd_sc_hd__and2_1 _5686_ (.A(net442),
    .B(net781),
    .X(_0842_));
 sky130_fd_sc_hd__and2_1 _5687_ (.A(net441),
    .B(net791),
    .X(_0843_));
 sky130_fd_sc_hd__or3b_2 _5688_ (.A(net2319),
    .B(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .C_N(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .X(_2726_));
 sky130_fd_sc_hd__nor2_4 _5689_ (.A(_1899_),
    .B(_2726_),
    .Y(_2727_));
 sky130_fd_sc_hd__or2_4 _5690_ (.A(_1899_),
    .B(_2726_),
    .X(_2728_));
 sky130_fd_sc_hd__nor2_2 _5691_ (.A(_1898_),
    .B(_1902_),
    .Y(_2729_));
 sky130_fd_sc_hd__or2_4 _5692_ (.A(_1898_),
    .B(_1902_),
    .X(_2730_));
 sky130_fd_sc_hd__nor2_2 _5693_ (.A(_2727_),
    .B(_2729_),
    .Y(_2731_));
 sky130_fd_sc_hd__nand2_4 _5694_ (.A(_2728_),
    .B(_2730_),
    .Y(_2732_));
 sky130_fd_sc_hd__mux4_1 _5695_ (.A0(_1654_),
    .A1(_1667_),
    .A2(_1700_),
    .A3(_1683_),
    .S0(net193),
    .S1(net189),
    .X(_2733_));
 sky130_fd_sc_hd__mux4_1 _5696_ (.A0(_1708_),
    .A1(_1724_),
    .A2(_1731_),
    .A3(_1742_),
    .S0(net189),
    .S1(net191),
    .X(_2734_));
 sky130_fd_sc_hd__mux2_1 _5697_ (.A0(_2733_),
    .A1(_2734_),
    .S(net197),
    .X(_2735_));
 sky130_fd_sc_hd__mux2_1 _5698_ (.A0(_1754_),
    .A1(_1778_),
    .S(net191),
    .X(_2736_));
 sky130_fd_sc_hd__mux4_1 _5699_ (.A0(_1754_),
    .A1(_1770_),
    .A2(_1778_),
    .A3(_1789_),
    .S0(net188),
    .S1(net191),
    .X(_2737_));
 sky130_fd_sc_hd__mux2_1 _5700_ (.A0(_1815_),
    .A1(_1834_),
    .S(net191),
    .X(_2738_));
 sky130_fd_sc_hd__mux2_1 _5701_ (.A0(_1802_),
    .A1(_1823_),
    .S(net190),
    .X(_2739_));
 sky130_fd_sc_hd__mux2_1 _5702_ (.A0(_2738_),
    .A1(_2739_),
    .S(net187),
    .X(_2740_));
 sky130_fd_sc_hd__mux2_1 _5703_ (.A0(_2737_),
    .A1(_2740_),
    .S(net197),
    .X(_2741_));
 sky130_fd_sc_hd__mux2_1 _5704_ (.A0(_2735_),
    .A1(_2741_),
    .S(net202),
    .X(_2742_));
 sky130_fd_sc_hd__mux2_1 _5705_ (.A0(_1513_),
    .A1(_1521_),
    .S(net190),
    .X(_2743_));
 sky130_fd_sc_hd__mux2_1 _5706_ (.A0(_1533_),
    .A1(_1545_),
    .S(net191),
    .X(_2744_));
 sky130_fd_sc_hd__mux2_1 _5707_ (.A0(_2743_),
    .A1(_2744_),
    .S(net186),
    .X(_2745_));
 sky130_fd_sc_hd__mux2_1 _5708_ (.A0(_1621_),
    .A1(_1640_),
    .S(_1681_),
    .X(_2746_));
 sky130_fd_sc_hd__mux2_1 _5709_ (.A0(_1605_),
    .A1(_1629_),
    .S(net191),
    .X(_2747_));
 sky130_fd_sc_hd__mux2_1 _5710_ (.A0(_2746_),
    .A1(_2747_),
    .S(net186),
    .X(_2748_));
 sky130_fd_sc_hd__mux2_1 _5711_ (.A0(_2745_),
    .A1(_2748_),
    .S(net194),
    .X(_2749_));
 sky130_fd_sc_hd__mux2_1 _5712_ (.A0(_1438_),
    .A1(_1487_),
    .S(net193),
    .X(_2750_));
 sky130_fd_sc_hd__mux2_1 _5713_ (.A0(_1471_),
    .A1(_1494_),
    .S(_1681_),
    .X(_2751_));
 sky130_fd_sc_hd__mux2_1 _5714_ (.A0(_2750_),
    .A1(_2751_),
    .S(net186),
    .X(_2752_));
 sky130_fd_sc_hd__mux2_1 _5715_ (.A0(_1572_),
    .A1(_1580_),
    .S(_1681_),
    .X(_2753_));
 sky130_fd_sc_hd__mux2_1 _5716_ (.A0(_1557_),
    .A1(_1594_),
    .S(_1681_),
    .X(_2754_));
 sky130_fd_sc_hd__mux2_1 _5717_ (.A0(_2753_),
    .A1(_2754_),
    .S(net186),
    .X(_2755_));
 sky130_fd_sc_hd__mux2_1 _5718_ (.A0(_2752_),
    .A1(_2755_),
    .S(net195),
    .X(_2756_));
 sky130_fd_sc_hd__mux2_2 _5719_ (.A0(_2749_),
    .A1(_2756_),
    .S(net202),
    .X(_2757_));
 sky130_fd_sc_hd__mux2_1 _5720_ (.A0(_2742_),
    .A1(_2757_),
    .S(net182),
    .X(_2758_));
 sky130_fd_sc_hd__inv_2 _5721_ (.A(_2758_),
    .Y(_2759_));
 sky130_fd_sc_hd__nor3_4 _5722_ (.A(net2340),
    .B(_1898_),
    .C(_1900_),
    .Y(_2760_));
 sky130_fd_sc_hd__or3_2 _5723_ (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .B(_1898_),
    .C(_1900_),
    .X(_2761_));
 sky130_fd_sc_hd__nor2_1 _5724_ (.A(net2358),
    .B(net2336),
    .Y(_2762_));
 sky130_fd_sc_hd__o31a_1 _5725_ (.A1(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .A2(net2336),
    .A3(_1897_),
    .B1(net354),
    .X(_2763_));
 sky130_fd_sc_hd__and2b_1 _5726_ (.A_N(_1902_),
    .B(_2762_),
    .X(_2764_));
 sky130_fd_sc_hd__or3_2 _5727_ (.A(net2358),
    .B(net2336),
    .C(_1902_),
    .X(_2765_));
 sky130_fd_sc_hd__nand2_1 _5728_ (.A(net302),
    .B(_2765_),
    .Y(_2766_));
 sky130_fd_sc_hd__nor2_1 _5729_ (.A(net2336),
    .B(_2726_),
    .Y(_2767_));
 sky130_fd_sc_hd__or2_1 _5730_ (.A(net2336),
    .B(_2726_),
    .X(_2768_));
 sky130_fd_sc_hd__nor2_1 _5731_ (.A(net2400),
    .B(_2768_),
    .Y(_2769_));
 sky130_fd_sc_hd__and4bb_2 _5732_ (.A_N(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ),
    .B_N(net2315),
    .C(net2340),
    .D(_2762_),
    .X(_2770_));
 sky130_fd_sc_hd__and4b_1 _5733_ (.A_N(net350),
    .B(_2731_),
    .C(_1903_),
    .D(_2768_),
    .X(_2771_));
 sky130_fd_sc_hd__and3_2 _5734_ (.A(net302),
    .B(_2765_),
    .C(_2771_),
    .X(_2772_));
 sky130_fd_sc_hd__a221o_1 _5735_ (.A1(_1686_),
    .A2(net300),
    .B1(net350),
    .B2(net191),
    .C1(net211),
    .X(_2773_));
 sky130_fd_sc_hd__a21oi_1 _5736_ (.A1(_1687_),
    .A2(_2766_),
    .B1(_2773_),
    .Y(_2774_));
 sky130_fd_sc_hd__and2_4 _5737_ (.A(net2358),
    .B(_2767_),
    .X(_2775_));
 sky130_fd_sc_hd__nand2_4 _5738_ (.A(net2358),
    .B(_2767_),
    .Y(_2776_));
 sky130_fd_sc_hd__nor2_4 _5739_ (.A(net182),
    .B(_2776_),
    .Y(_2777_));
 sky130_fd_sc_hd__nand2_2 _5740_ (.A(_1721_),
    .B(_2775_),
    .Y(_2778_));
 sky130_fd_sc_hd__o41a_1 _5741_ (.A1(net202),
    .A2(net197),
    .A3(_1846_),
    .A4(_2778_),
    .B1(_2774_),
    .X(_2779_));
 sky130_fd_sc_hd__o221a_1 _5742_ (.A1(_1894_),
    .A2(net2341),
    .B1(_2731_),
    .B2(_2759_),
    .C1(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__a211oi_1 _5743_ (.A1(_1685_),
    .A2(net211),
    .B1(net2342),
    .C1(net466),
    .Y(_0844_));
 sky130_fd_sc_hd__mux2_1 _5744_ (.A0(_1521_),
    .A1(_1533_),
    .S(net190),
    .X(_2781_));
 sky130_fd_sc_hd__mux4_1 _5745_ (.A0(_1521_),
    .A1(_1533_),
    .A2(_1545_),
    .A3(_1621_),
    .S0(net190),
    .S1(net185),
    .X(_2782_));
 sky130_fd_sc_hd__mux4_1 _5746_ (.A0(_1487_),
    .A1(_1605_),
    .A2(_1629_),
    .A3(_1640_),
    .S0(net188),
    .S1(_1680_),
    .X(_2783_));
 sky130_fd_sc_hd__mux2_1 _5747_ (.A0(_2782_),
    .A1(_2783_),
    .S(net195),
    .X(_2784_));
 sky130_fd_sc_hd__nor2_1 _5748_ (.A(net203),
    .B(_2784_),
    .Y(_2785_));
 sky130_fd_sc_hd__mux4_1 _5749_ (.A0(_1438_),
    .A1(_1471_),
    .A2(_1494_),
    .A3(_1572_),
    .S0(_1681_),
    .S1(net186),
    .X(_2786_));
 sky130_fd_sc_hd__nor2_1 _5750_ (.A(net195),
    .B(_2786_),
    .Y(_2787_));
 sky130_fd_sc_hd__mux2_1 _5751_ (.A0(_1557_),
    .A1(_1580_),
    .S(net193),
    .X(_2788_));
 sky130_fd_sc_hd__and2_1 _5752_ (.A(net189),
    .B(_2788_),
    .X(_2789_));
 sky130_fd_sc_hd__a21oi_1 _5753_ (.A1(_1594_),
    .A2(net186),
    .B1(_2789_),
    .Y(_2790_));
 sky130_fd_sc_hd__a21oi_1 _5754_ (.A1(net195),
    .A2(_2790_),
    .B1(_2787_),
    .Y(_2791_));
 sky130_fd_sc_hd__o21ba_1 _5755_ (.A1(net205),
    .A2(_2791_),
    .B1_N(_2785_),
    .X(_2792_));
 sky130_fd_sc_hd__nand2_1 _5756_ (.A(_1594_),
    .B(net193),
    .Y(_2793_));
 sky130_fd_sc_hd__o21ba_1 _5757_ (.A1(net189),
    .A2(_2793_),
    .B1_N(_2789_),
    .X(_2794_));
 sky130_fd_sc_hd__a21o_1 _5758_ (.A1(net195),
    .A2(_2794_),
    .B1(_2787_),
    .X(_2795_));
 sky130_fd_sc_hd__inv_2 _5759_ (.A(_2795_),
    .Y(_2796_));
 sky130_fd_sc_hd__a21oi_1 _5760_ (.A1(net203),
    .A2(_2795_),
    .B1(_2785_),
    .Y(_2797_));
 sky130_fd_sc_hd__a22o_1 _5761_ (.A1(_2727_),
    .A2(_2792_),
    .B1(_2797_),
    .B2(_2729_),
    .X(_2798_));
 sky130_fd_sc_hd__nand2_1 _5762_ (.A(net181),
    .B(_2798_),
    .Y(_2799_));
 sky130_fd_sc_hd__or3_1 _5763_ (.A(_1694_),
    .B(_1696_),
    .C(net355),
    .X(_2800_));
 sky130_fd_sc_hd__o21ai_1 _5764_ (.A1(_1694_),
    .A2(_1696_),
    .B1(net355),
    .Y(_2801_));
 sky130_fd_sc_hd__and3_1 _5765_ (.A(_1700_),
    .B(_2800_),
    .C(_2801_),
    .X(_2802_));
 sky130_fd_sc_hd__a21o_1 _5766_ (.A1(_2800_),
    .A2(_2801_),
    .B1(_1700_),
    .X(_2803_));
 sky130_fd_sc_hd__and2b_1 _5767_ (.A_N(_2802_),
    .B(_2803_),
    .X(_2804_));
 sky130_fd_sc_hd__mux2_1 _5768_ (.A0(_1683_),
    .A1(net355),
    .S(net193),
    .X(_2805_));
 sky130_fd_sc_hd__xnor2_1 _5769_ (.A(_2804_),
    .B(_2805_),
    .Y(_2806_));
 sky130_fd_sc_hd__a221o_1 _5770_ (.A1(_1702_),
    .A2(net300),
    .B1(net350),
    .B2(net187),
    .C1(net211),
    .X(_2807_));
 sky130_fd_sc_hd__a21oi_1 _5771_ (.A1(net352),
    .A2(_2804_),
    .B1(_2807_),
    .Y(_2808_));
 sky130_fd_sc_hd__mux2_1 _5772_ (.A0(_1684_),
    .A1(_1701_),
    .S(net193),
    .X(_2809_));
 sky130_fd_sc_hd__or3_1 _5773_ (.A(net196),
    .B(net187),
    .C(_2809_),
    .X(_2810_));
 sky130_fd_sc_hd__or2_1 _5774_ (.A(net201),
    .B(_2810_),
    .X(_2811_));
 sky130_fd_sc_hd__o221a_1 _5775_ (.A1(net302),
    .A2(_2806_),
    .B1(_2811_),
    .B2(_2778_),
    .C1(_2808_),
    .X(_2812_));
 sky130_fd_sc_hd__mux4_1 _5776_ (.A0(_1654_),
    .A1(_1700_),
    .A2(_1724_),
    .A3(_1667_),
    .S0(net189),
    .S1(net191),
    .X(_2813_));
 sky130_fd_sc_hd__mux4_1 _5777_ (.A0(_1708_),
    .A1(_1742_),
    .A2(_1770_),
    .A3(_1731_),
    .S0(net192),
    .S1(net187),
    .X(_2814_));
 sky130_fd_sc_hd__mux2_1 _5778_ (.A0(_2813_),
    .A1(_2814_),
    .S(net196),
    .X(_2815_));
 sky130_fd_sc_hd__mux2_1 _5779_ (.A0(_1778_),
    .A1(_1815_),
    .S(net191),
    .X(_2816_));
 sky130_fd_sc_hd__mux4_1 _5780_ (.A0(_1754_),
    .A1(_1789_),
    .A2(_1815_),
    .A3(_1778_),
    .S0(net193),
    .S1(net187),
    .X(_2817_));
 sky130_fd_sc_hd__mux2_1 _5781_ (.A0(_1513_),
    .A1(_1823_),
    .S(net192),
    .X(_2818_));
 sky130_fd_sc_hd__mux2_1 _5782_ (.A0(_1802_),
    .A1(_1834_),
    .S(net192),
    .X(_2819_));
 sky130_fd_sc_hd__mux2_1 _5783_ (.A0(_2818_),
    .A1(_2819_),
    .S(net188),
    .X(_2820_));
 sky130_fd_sc_hd__mux2_1 _5784_ (.A0(_2817_),
    .A1(_2820_),
    .S(net196),
    .X(_2821_));
 sky130_fd_sc_hd__mux2_1 _5785_ (.A0(_2815_),
    .A1(_2821_),
    .S(net201),
    .X(_2822_));
 sky130_fd_sc_hd__or3b_1 _5786_ (.A(net181),
    .B(_2731_),
    .C_N(_2822_),
    .X(_2823_));
 sky130_fd_sc_hd__a32o_1 _5787_ (.A1(_2799_),
    .A2(_2812_),
    .A3(_2823_),
    .B1(net211),
    .B2(_1703_),
    .X(_2824_));
 sky130_fd_sc_hd__nor2_1 _5788_ (.A(net467),
    .B(net2395),
    .Y(_0845_));
 sky130_fd_sc_hd__mux2_1 _5789_ (.A0(_1667_),
    .A1(_1700_),
    .S(net191),
    .X(_2825_));
 sky130_fd_sc_hd__o21bai_1 _5790_ (.A1(net186),
    .A2(_2825_),
    .B1_N(_1845_),
    .Y(_2826_));
 sky130_fd_sc_hd__inv_2 _5791_ (.A(_2826_),
    .Y(_2827_));
 sky130_fd_sc_hd__nor2_1 _5792_ (.A(net197),
    .B(_2826_),
    .Y(_2828_));
 sky130_fd_sc_hd__nor2_2 _5793_ (.A(net202),
    .B(_2776_),
    .Y(_2829_));
 sky130_fd_sc_hd__mux4_1 _5794_ (.A0(_1654_),
    .A1(_1667_),
    .A2(_1742_),
    .A3(_1724_),
    .S0(net193),
    .S1(net187),
    .X(_2830_));
 sky130_fd_sc_hd__mux4_1 _5795_ (.A0(_1708_),
    .A1(_1731_),
    .A2(_1770_),
    .A3(_1789_),
    .S0(net190),
    .S1(net187),
    .X(_2831_));
 sky130_fd_sc_hd__mux2_1 _5796_ (.A0(_2830_),
    .A1(_2831_),
    .S(net196),
    .X(_2832_));
 sky130_fd_sc_hd__mux2_1 _5797_ (.A0(_2736_),
    .A1(_2738_),
    .S(net187),
    .X(_2833_));
 sky130_fd_sc_hd__mux2_1 _5798_ (.A0(_2739_),
    .A1(_2743_),
    .S(net185),
    .X(_2834_));
 sky130_fd_sc_hd__mux2_1 _5799_ (.A0(_2833_),
    .A1(_2834_),
    .S(net196),
    .X(_2835_));
 sky130_fd_sc_hd__mux2_1 _5800_ (.A0(_2832_),
    .A1(_2835_),
    .S(net201),
    .X(_2836_));
 sky130_fd_sc_hd__a22o_1 _5801_ (.A1(_2828_),
    .A2(_2829_),
    .B1(_2836_),
    .B2(_2732_),
    .X(_2837_));
 sky130_fd_sc_hd__mux2_1 _5802_ (.A0(_2751_),
    .A1(_2753_),
    .S(net186),
    .X(_2838_));
 sky130_fd_sc_hd__nor2_1 _5803_ (.A(net194),
    .B(_2838_),
    .Y(_2839_));
 sky130_fd_sc_hd__nand2_1 _5804_ (.A(net189),
    .B(_2754_),
    .Y(_2840_));
 sky130_fd_sc_hd__a21oi_1 _5805_ (.A1(net194),
    .A2(_2840_),
    .B1(_2839_),
    .Y(_2841_));
 sky130_fd_sc_hd__nor2_1 _5806_ (.A(net204),
    .B(_2841_),
    .Y(_2842_));
 sky130_fd_sc_hd__mux2_1 _5807_ (.A0(_2744_),
    .A1(_2746_),
    .S(net186),
    .X(_2843_));
 sky130_fd_sc_hd__mux2_1 _5808_ (.A0(_2747_),
    .A1(_2750_),
    .S(net186),
    .X(_2844_));
 sky130_fd_sc_hd__mux2_1 _5809_ (.A0(_2843_),
    .A1(_2844_),
    .S(net194),
    .X(_2845_));
 sky130_fd_sc_hd__nor2_1 _5810_ (.A(net203),
    .B(_2845_),
    .Y(_2846_));
 sky130_fd_sc_hd__or3_1 _5811_ (.A(_2730_),
    .B(_2842_),
    .C(_2846_),
    .X(_2847_));
 sky130_fd_sc_hd__o21a_1 _5812_ (.A1(_1595_),
    .A2(net189),
    .B1(_2840_),
    .X(_2848_));
 sky130_fd_sc_hd__a21oi_1 _5813_ (.A1(net194),
    .A2(_2848_),
    .B1(_2839_),
    .Y(_2849_));
 sky130_fd_sc_hd__nor2_1 _5814_ (.A(net204),
    .B(_2849_),
    .Y(_2850_));
 sky130_fd_sc_hd__or3_1 _5815_ (.A(_2728_),
    .B(_2846_),
    .C(_2850_),
    .X(_2851_));
 sky130_fd_sc_hd__a21oi_1 _5816_ (.A1(_2847_),
    .A2(_2851_),
    .B1(net183),
    .Y(_2852_));
 sky130_fd_sc_hd__o21a_1 _5817_ (.A1(_2802_),
    .A2(_2805_),
    .B1(_2803_),
    .X(_2853_));
 sky130_fd_sc_hd__nand2_1 _5818_ (.A(net199),
    .B(net354),
    .Y(_2854_));
 sky130_fd_sc_hd__nand2_1 _5819_ (.A(net196),
    .B(net355),
    .Y(_2855_));
 sky130_fd_sc_hd__and3_1 _5820_ (.A(_1667_),
    .B(_2854_),
    .C(_2855_),
    .X(_2856_));
 sky130_fd_sc_hd__a21o_1 _5821_ (.A1(_2854_),
    .A2(_2855_),
    .B1(_1667_),
    .X(_2857_));
 sky130_fd_sc_hd__and2b_1 _5822_ (.A_N(_2856_),
    .B(_2857_),
    .X(_2858_));
 sky130_fd_sc_hd__xnor2_1 _5823_ (.A(_2853_),
    .B(_2858_),
    .Y(_2859_));
 sky130_fd_sc_hd__o21a_1 _5824_ (.A1(_1667_),
    .A2(net196),
    .B1(net300),
    .X(_2860_));
 sky130_fd_sc_hd__a211o_1 _5825_ (.A1(net196),
    .A2(net350),
    .B1(net210),
    .C1(_2860_),
    .X(_2861_));
 sky130_fd_sc_hd__o22ai_1 _5826_ (.A1(_1673_),
    .A2(_2765_),
    .B1(_2859_),
    .B2(net302),
    .Y(_2862_));
 sky130_fd_sc_hd__a211o_1 _5827_ (.A1(net184),
    .A2(_2837_),
    .B1(_2861_),
    .C1(_2862_),
    .X(_2863_));
 sky130_fd_sc_hd__a21bo_1 _5828_ (.A1(_1667_),
    .A2(net196),
    .B1_N(net210),
    .X(_2864_));
 sky130_fd_sc_hd__o211a_1 _5829_ (.A1(_2852_),
    .A2(_2863_),
    .B1(_2864_),
    .C1(net459),
    .X(_0846_));
 sky130_fd_sc_hd__mux4_1 _5830_ (.A0(_1545_),
    .A1(_1621_),
    .A2(_1640_),
    .A3(_1605_),
    .S0(net190),
    .S1(net185),
    .X(_2865_));
 sky130_fd_sc_hd__mux4_1 _5831_ (.A0(_1438_),
    .A1(_1471_),
    .A2(_1629_),
    .A3(_1487_),
    .S0(net190),
    .S1(net188),
    .X(_2866_));
 sky130_fd_sc_hd__mux2_1 _5832_ (.A0(_2865_),
    .A1(_2866_),
    .S(net195),
    .X(_2867_));
 sky130_fd_sc_hd__mux4_1 _5833_ (.A0(_1494_),
    .A1(_1572_),
    .A2(_1580_),
    .A3(_1557_),
    .S0(net190),
    .S1(net185),
    .X(_2868_));
 sky130_fd_sc_hd__nand2_1 _5834_ (.A(net198),
    .B(_2868_),
    .Y(_2869_));
 sky130_fd_sc_hd__nand2_1 _5835_ (.A(_1594_),
    .B(net194),
    .Y(_2870_));
 sky130_fd_sc_hd__nand2_1 _5836_ (.A(_2869_),
    .B(_2870_),
    .Y(_2871_));
 sky130_fd_sc_hd__mux2_1 _5837_ (.A0(_2867_),
    .A1(_2871_),
    .S(net203),
    .X(_2872_));
 sky130_fd_sc_hd__or2_1 _5838_ (.A(net186),
    .B(_2793_),
    .X(_2873_));
 sky130_fd_sc_hd__o21a_1 _5839_ (.A1(net200),
    .A2(_2873_),
    .B1(_2869_),
    .X(_2874_));
 sky130_fd_sc_hd__inv_2 _5840_ (.A(_2874_),
    .Y(_2875_));
 sky130_fd_sc_hd__mux2_1 _5841_ (.A0(_2867_),
    .A1(_2875_),
    .S(net203),
    .X(_2876_));
 sky130_fd_sc_hd__a22o_1 _5842_ (.A1(_2727_),
    .A2(_2872_),
    .B1(_2876_),
    .B2(_2729_),
    .X(_2877_));
 sky130_fd_sc_hd__xnor2_1 _5843_ (.A(net206),
    .B(net355),
    .Y(_2878_));
 sky130_fd_sc_hd__and2_1 _5844_ (.A(_1654_),
    .B(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__nand2_1 _5845_ (.A(_1654_),
    .B(_2878_),
    .Y(_2880_));
 sky130_fd_sc_hd__nor2_1 _5846_ (.A(_1654_),
    .B(_2878_),
    .Y(_2881_));
 sky130_fd_sc_hd__nor2_1 _5847_ (.A(_2879_),
    .B(_2881_),
    .Y(_2882_));
 sky130_fd_sc_hd__o21ai_1 _5848_ (.A1(_2853_),
    .A2(_2856_),
    .B1(_2857_),
    .Y(_2883_));
 sky130_fd_sc_hd__nand2_1 _5849_ (.A(_2882_),
    .B(_2883_),
    .Y(_2884_));
 sky130_fd_sc_hd__or2_1 _5850_ (.A(_2882_),
    .B(_2883_),
    .X(_2885_));
 sky130_fd_sc_hd__a21oi_1 _5851_ (.A1(_2884_),
    .A2(_2885_),
    .B1(net302),
    .Y(_2886_));
 sky130_fd_sc_hd__mux4_2 _5852_ (.A0(_1654_),
    .A1(_1667_),
    .A2(_1700_),
    .A3(_1683_),
    .S0(net191),
    .S1(net186),
    .X(_2887_));
 sky130_fd_sc_hd__and3_1 _5853_ (.A(net206),
    .B(net199),
    .C(_2887_),
    .X(_2888_));
 sky130_fd_sc_hd__a221o_1 _5854_ (.A1(_1661_),
    .A2(net300),
    .B1(net350),
    .B2(net201),
    .C1(net210),
    .X(_2889_));
 sky130_fd_sc_hd__a22o_1 _5855_ (.A1(net352),
    .A2(_2882_),
    .B1(_2888_),
    .B2(_2777_),
    .X(_2890_));
 sky130_fd_sc_hd__mux4_1 _5856_ (.A0(_1654_),
    .A1(_1724_),
    .A2(_1742_),
    .A3(_1708_),
    .S0(net190),
    .S1(net185),
    .X(_2891_));
 sky130_fd_sc_hd__mux4_1 _5857_ (.A0(_1731_),
    .A1(_1770_),
    .A2(_1789_),
    .A3(_1754_),
    .S0(net190),
    .S1(net185),
    .X(_2892_));
 sky130_fd_sc_hd__mux2_1 _5858_ (.A0(_2891_),
    .A1(_2892_),
    .S(net196),
    .X(_2893_));
 sky130_fd_sc_hd__mux2_1 _5859_ (.A0(_2816_),
    .A1(_2819_),
    .S(net185),
    .X(_2894_));
 sky130_fd_sc_hd__mux2_1 _5860_ (.A0(_2781_),
    .A1(_2818_),
    .S(net188),
    .X(_2895_));
 sky130_fd_sc_hd__mux2_1 _5861_ (.A0(_2894_),
    .A1(_2895_),
    .S(net196),
    .X(_2896_));
 sky130_fd_sc_hd__mux2_1 _5862_ (.A0(_2893_),
    .A1(_2896_),
    .S(net201),
    .X(_2897_));
 sky130_fd_sc_hd__a311o_1 _5863_ (.A1(net184),
    .A2(_2732_),
    .A3(_2897_),
    .B1(_2890_),
    .C1(_2889_),
    .X(_2898_));
 sky130_fd_sc_hd__a211oi_1 _5864_ (.A1(net181),
    .A2(_2877_),
    .B1(_2886_),
    .C1(_2898_),
    .Y(_2899_));
 sky130_fd_sc_hd__a211oi_1 _5865_ (.A1(_1660_),
    .A2(net210),
    .B1(_2899_),
    .C1(net466),
    .Y(_0847_));
 sky130_fd_sc_hd__a21o_1 _5866_ (.A1(_2880_),
    .A2(_2883_),
    .B1(_2881_),
    .X(_2900_));
 sky130_fd_sc_hd__xnor2_1 _5867_ (.A(net184),
    .B(net355),
    .Y(_2901_));
 sky130_fd_sc_hd__nand2_1 _5868_ (.A(_1724_),
    .B(_2901_),
    .Y(_2902_));
 sky130_fd_sc_hd__nor2_1 _5869_ (.A(_1724_),
    .B(_2901_),
    .Y(_2903_));
 sky130_fd_sc_hd__or2_1 _5870_ (.A(_1724_),
    .B(_2901_),
    .X(_2904_));
 sky130_fd_sc_hd__nand2_1 _5871_ (.A(_2902_),
    .B(_2904_),
    .Y(_2905_));
 sky130_fd_sc_hd__xnor2_1 _5872_ (.A(_2900_),
    .B(_2905_),
    .Y(_2906_));
 sky130_fd_sc_hd__mux2_1 _5873_ (.A0(_2748_),
    .A1(_2752_),
    .S(net195),
    .X(_2907_));
 sky130_fd_sc_hd__and2_1 _5874_ (.A(net200),
    .B(_2755_),
    .X(_2908_));
 sky130_fd_sc_hd__a21o_1 _5875_ (.A1(_1594_),
    .A2(net194),
    .B1(_2908_),
    .X(_2909_));
 sky130_fd_sc_hd__mux2_1 _5876_ (.A0(_2907_),
    .A1(_2909_),
    .S(net203),
    .X(_2910_));
 sky130_fd_sc_hd__mux4_1 _5877_ (.A0(_1654_),
    .A1(_1700_),
    .A2(_1724_),
    .A3(_1667_),
    .S0(net187),
    .S1(net193),
    .X(_2911_));
 sky130_fd_sc_hd__mux2_1 _5878_ (.A0(_1847_),
    .A1(_2911_),
    .S(net200),
    .X(_2912_));
 sky130_fd_sc_hd__mux2_1 _5879_ (.A0(_2734_),
    .A1(_2737_),
    .S(net197),
    .X(_2913_));
 sky130_fd_sc_hd__mux2_1 _5880_ (.A0(_2740_),
    .A1(_2745_),
    .S(net194),
    .X(_2914_));
 sky130_fd_sc_hd__or4_1 _5881_ (.A(net204),
    .B(_1721_),
    .C(_2727_),
    .D(_2908_),
    .X(_2915_));
 sky130_fd_sc_hd__mux4_1 _5882_ (.A0(_2907_),
    .A1(_2909_),
    .A2(_2913_),
    .A3(_2914_),
    .S0(net202),
    .S1(net184),
    .X(_2916_));
 sky130_fd_sc_hd__a221o_1 _5883_ (.A1(_1725_),
    .A2(net300),
    .B1(net350),
    .B2(net182),
    .C1(net211),
    .X(_2917_));
 sky130_fd_sc_hd__a31o_1 _5884_ (.A1(_1725_),
    .A2(_1726_),
    .A3(net352),
    .B1(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__a31o_1 _5885_ (.A1(net207),
    .A2(_2777_),
    .A3(_2912_),
    .B1(_2918_),
    .X(_2919_));
 sky130_fd_sc_hd__a31o_1 _5886_ (.A1(_2732_),
    .A2(_2915_),
    .A3(_2916_),
    .B1(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__o21ba_1 _5887_ (.A1(net302),
    .A2(_2906_),
    .B1_N(_2920_),
    .X(_2921_));
 sky130_fd_sc_hd__a211oi_2 _5888_ (.A1(_1726_),
    .A2(net211),
    .B1(_2921_),
    .C1(net468),
    .Y(_0848_));
 sky130_fd_sc_hd__xnor2_1 _5889_ (.A(_1745_),
    .B(net354),
    .Y(_2922_));
 sky130_fd_sc_hd__and2_1 _5890_ (.A(_1742_),
    .B(_2922_),
    .X(_2923_));
 sky130_fd_sc_hd__nand2_1 _5891_ (.A(_1742_),
    .B(_2922_),
    .Y(_2924_));
 sky130_fd_sc_hd__nor2_1 _5892_ (.A(_1742_),
    .B(_2922_),
    .Y(_2925_));
 sky130_fd_sc_hd__nor2_1 _5893_ (.A(_2923_),
    .B(_2925_),
    .Y(_2926_));
 sky130_fd_sc_hd__a21o_1 _5894_ (.A1(_2900_),
    .A2(_2902_),
    .B1(_2903_),
    .X(_2927_));
 sky130_fd_sc_hd__xor2_1 _5895_ (.A(_2926_),
    .B(_2927_),
    .X(_2928_));
 sky130_fd_sc_hd__mux2_1 _5896_ (.A0(_2783_),
    .A1(_2786_),
    .S(net195),
    .X(_2929_));
 sky130_fd_sc_hd__nor2_1 _5897_ (.A(net203),
    .B(_2929_),
    .Y(_2930_));
 sky130_fd_sc_hd__nor2_1 _5898_ (.A(net194),
    .B(_2794_),
    .Y(_2931_));
 sky130_fd_sc_hd__nor2_1 _5899_ (.A(net205),
    .B(_2931_),
    .Y(_2932_));
 sky130_fd_sc_hd__or3_1 _5900_ (.A(_2730_),
    .B(_2930_),
    .C(_2932_),
    .X(_2933_));
 sky130_fd_sc_hd__o21a_1 _5901_ (.A1(net194),
    .A2(_2790_),
    .B1(_2870_),
    .X(_2934_));
 sky130_fd_sc_hd__a21oi_1 _5902_ (.A1(net203),
    .A2(_2934_),
    .B1(_2930_),
    .Y(_2935_));
 sky130_fd_sc_hd__a21bo_1 _5903_ (.A1(_2727_),
    .A2(_2935_),
    .B1_N(_2933_),
    .X(_2936_));
 sky130_fd_sc_hd__a221o_1 _5904_ (.A1(_1746_),
    .A2(net300),
    .B1(net350),
    .B2(_1745_),
    .C1(net211),
    .X(_2937_));
 sky130_fd_sc_hd__mux4_1 _5905_ (.A0(_1654_),
    .A1(_1667_),
    .A2(_1742_),
    .A3(_1724_),
    .S0(net190),
    .S1(net188),
    .X(_2938_));
 sky130_fd_sc_hd__nand2_1 _5906_ (.A(net199),
    .B(_2938_),
    .Y(_2939_));
 sky130_fd_sc_hd__o31a_1 _5907_ (.A1(net199),
    .A2(net187),
    .A3(_2809_),
    .B1(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__mux2_1 _5908_ (.A0(_2814_),
    .A1(_2817_),
    .S(net196),
    .X(_2941_));
 sky130_fd_sc_hd__mux2_1 _5909_ (.A0(_2782_),
    .A1(_2820_),
    .S(net199),
    .X(_2942_));
 sky130_fd_sc_hd__mux2_1 _5910_ (.A0(_2941_),
    .A1(_2942_),
    .S(net201),
    .X(_2943_));
 sky130_fd_sc_hd__inv_2 _5911_ (.A(_2943_),
    .Y(_2944_));
 sky130_fd_sc_hd__o32a_1 _5912_ (.A1(net201),
    .A2(_2776_),
    .A3(_2940_),
    .B1(_2944_),
    .B2(_2731_),
    .X(_2945_));
 sky130_fd_sc_hd__a22o_1 _5913_ (.A1(net352),
    .A2(_2926_),
    .B1(_2936_),
    .B2(net181),
    .X(_2946_));
 sky130_fd_sc_hd__nor2_1 _5914_ (.A(_2937_),
    .B(_2946_),
    .Y(_2947_));
 sky130_fd_sc_hd__o22a_1 _5915_ (.A1(net302),
    .A2(_2928_),
    .B1(_2945_),
    .B2(net181),
    .X(_2948_));
 sky130_fd_sc_hd__a221oi_4 _5916_ (.A1(net2389),
    .A2(net211),
    .B1(_2947_),
    .B2(_2948_),
    .C1(net467),
    .Y(_0849_));
 sky130_fd_sc_hd__a21o_1 _5917_ (.A1(_2924_),
    .A2(_2927_),
    .B1(_2925_),
    .X(_2949_));
 sky130_fd_sc_hd__xnor2_1 _5918_ (.A(_1711_),
    .B(net354),
    .Y(_2950_));
 sky130_fd_sc_hd__nand2_1 _5919_ (.A(_1708_),
    .B(_2950_),
    .Y(_2951_));
 sky130_fd_sc_hd__nor2_1 _5920_ (.A(_1708_),
    .B(_2950_),
    .Y(_2952_));
 sky130_fd_sc_hd__or2_1 _5921_ (.A(_1708_),
    .B(_2950_),
    .X(_2953_));
 sky130_fd_sc_hd__nand2_1 _5922_ (.A(_2951_),
    .B(_2953_),
    .Y(_2954_));
 sky130_fd_sc_hd__xnor2_1 _5923_ (.A(_2949_),
    .B(_2954_),
    .Y(_2955_));
 sky130_fd_sc_hd__mux2_1 _5924_ (.A0(_2838_),
    .A1(_2844_),
    .S(net200),
    .X(_2956_));
 sky130_fd_sc_hd__or2_1 _5925_ (.A(net203),
    .B(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__nor2_1 _5926_ (.A(net194),
    .B(_2840_),
    .Y(_2958_));
 sky130_fd_sc_hd__o211a_1 _5927_ (.A1(net204),
    .A2(_2958_),
    .B1(_2957_),
    .C1(_2729_),
    .X(_2959_));
 sky130_fd_sc_hd__o21ai_1 _5928_ (.A1(net194),
    .A2(_2848_),
    .B1(_2870_),
    .Y(_2960_));
 sky130_fd_sc_hd__o21ai_1 _5929_ (.A1(net204),
    .A2(_2960_),
    .B1(_2957_),
    .Y(_2961_));
 sky130_fd_sc_hd__nor2_1 _5930_ (.A(_2728_),
    .B(_2961_),
    .Y(_2962_));
 sky130_fd_sc_hd__o21a_1 _5931_ (.A1(_2959_),
    .A2(_2962_),
    .B1(net182),
    .X(_2963_));
 sky130_fd_sc_hd__a221o_1 _5932_ (.A1(_1712_),
    .A2(net300),
    .B1(net350),
    .B2(_1711_),
    .C1(net211),
    .X(_2964_));
 sky130_fd_sc_hd__a211oi_1 _5933_ (.A1(_1714_),
    .A2(net352),
    .B1(_2963_),
    .C1(_2964_),
    .Y(_2965_));
 sky130_fd_sc_hd__mux4_1 _5934_ (.A0(_1654_),
    .A1(_1724_),
    .A2(_1742_),
    .A3(_1708_),
    .S0(net193),
    .S1(net189),
    .X(_2966_));
 sky130_fd_sc_hd__mux2_1 _5935_ (.A0(_2827_),
    .A1(_2966_),
    .S(net199),
    .X(_2967_));
 sky130_fd_sc_hd__nand2_1 _5936_ (.A(net207),
    .B(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__mux2_1 _5937_ (.A0(_2831_),
    .A1(_2833_),
    .S(net196),
    .X(_2969_));
 sky130_fd_sc_hd__mux2_1 _5938_ (.A0(_2834_),
    .A1(_2843_),
    .S(net194),
    .X(_2970_));
 sky130_fd_sc_hd__mux2_1 _5939_ (.A0(_2969_),
    .A1(_2970_),
    .S(net202),
    .X(_2971_));
 sky130_fd_sc_hd__o2bb2a_1 _5940_ (.A1_N(_2732_),
    .A2_N(_2971_),
    .B1(_2968_),
    .B2(_2776_),
    .X(_2972_));
 sky130_fd_sc_hd__o22a_1 _5941_ (.A1(net302),
    .A2(_2955_),
    .B1(_2972_),
    .B2(net181),
    .X(_2973_));
 sky130_fd_sc_hd__a221oi_2 _5942_ (.A1(_1713_),
    .A2(net211),
    .B1(_2965_),
    .B2(_2973_),
    .C1(net467),
    .Y(_0850_));
 sky130_fd_sc_hd__xnor2_1 _5943_ (.A(_1734_),
    .B(net354),
    .Y(_2974_));
 sky130_fd_sc_hd__and2_1 _5944_ (.A(_1731_),
    .B(_2974_),
    .X(_2975_));
 sky130_fd_sc_hd__nand2_1 _5945_ (.A(_1731_),
    .B(_2974_),
    .Y(_2976_));
 sky130_fd_sc_hd__nor2_1 _5946_ (.A(_1731_),
    .B(_2974_),
    .Y(_2977_));
 sky130_fd_sc_hd__nor2_1 _5947_ (.A(_2975_),
    .B(_2977_),
    .Y(_2978_));
 sky130_fd_sc_hd__a21o_1 _5948_ (.A1(_2949_),
    .A2(_2951_),
    .B1(_2952_),
    .X(_2979_));
 sky130_fd_sc_hd__xor2_1 _5949_ (.A(_2978_),
    .B(_2979_),
    .X(_2980_));
 sky130_fd_sc_hd__mux2_1 _5950_ (.A0(_2866_),
    .A1(_2868_),
    .S(net195),
    .X(_2981_));
 sky130_fd_sc_hd__nand2_1 _5951_ (.A(net205),
    .B(_2981_),
    .Y(_2982_));
 sky130_fd_sc_hd__nor2_1 _5952_ (.A(net194),
    .B(_2873_),
    .Y(_2983_));
 sky130_fd_sc_hd__nand2_1 _5953_ (.A(net203),
    .B(_2983_),
    .Y(_2984_));
 sky130_fd_sc_hd__a21oi_1 _5954_ (.A1(_2982_),
    .A2(_2984_),
    .B1(_2730_),
    .Y(_2985_));
 sky130_fd_sc_hd__nor2_2 _5955_ (.A(_1595_),
    .B(net204),
    .Y(_2986_));
 sky130_fd_sc_hd__nand2_1 _5956_ (.A(_1594_),
    .B(net203),
    .Y(_2987_));
 sky130_fd_sc_hd__nand2_1 _5957_ (.A(_2982_),
    .B(_2987_),
    .Y(_2988_));
 sky130_fd_sc_hd__a21o_1 _5958_ (.A1(_2727_),
    .A2(_2988_),
    .B1(_2985_),
    .X(_2989_));
 sky130_fd_sc_hd__a221o_1 _5959_ (.A1(_1735_),
    .A2(net300),
    .B1(net350),
    .B2(_1734_),
    .C1(net210),
    .X(_2990_));
 sky130_fd_sc_hd__a22o_1 _5960_ (.A1(net352),
    .A2(_2978_),
    .B1(_2989_),
    .B2(net182),
    .X(_2991_));
 sky130_fd_sc_hd__mux4_1 _5961_ (.A0(_1708_),
    .A1(_1724_),
    .A2(_1731_),
    .A3(_1742_),
    .S0(net185),
    .S1(net192),
    .X(_2992_));
 sky130_fd_sc_hd__mux2_1 _5962_ (.A0(_2887_),
    .A1(_2992_),
    .S(net199),
    .X(_2993_));
 sky130_fd_sc_hd__mux2_1 _5963_ (.A0(_2892_),
    .A1(_2894_),
    .S(net196),
    .X(_2994_));
 sky130_fd_sc_hd__mux2_1 _5964_ (.A0(_2865_),
    .A1(_2895_),
    .S(net198),
    .X(_2995_));
 sky130_fd_sc_hd__mux2_1 _5965_ (.A0(_2994_),
    .A1(_2995_),
    .S(net202),
    .X(_2996_));
 sky130_fd_sc_hd__a22o_1 _5966_ (.A1(_2829_),
    .A2(_2993_),
    .B1(_2996_),
    .B2(_2732_),
    .X(_2997_));
 sky130_fd_sc_hd__a2bb2o_1 _5967_ (.A1_N(net302),
    .A2_N(_2980_),
    .B1(_2997_),
    .B2(net184),
    .X(_2998_));
 sky130_fd_sc_hd__a21oi_1 _5968_ (.A1(_1736_),
    .A2(net210),
    .B1(net468),
    .Y(_2999_));
 sky130_fd_sc_hd__o31a_1 _5969_ (.A1(_2990_),
    .A2(_2991_),
    .A3(_2998_),
    .B1(_2999_),
    .X(_0851_));
 sky130_fd_sc_hd__a21o_1 _5970_ (.A1(_2976_),
    .A2(_2979_),
    .B1(_2977_),
    .X(_3000_));
 sky130_fd_sc_hd__xnor2_1 _5971_ (.A(_1767_),
    .B(net355),
    .Y(_3001_));
 sky130_fd_sc_hd__nand2_1 _5972_ (.A(_1770_),
    .B(_3001_),
    .Y(_3002_));
 sky130_fd_sc_hd__nor2_1 _5973_ (.A(_1770_),
    .B(_3001_),
    .Y(_3003_));
 sky130_fd_sc_hd__or2_1 _5974_ (.A(_1770_),
    .B(_3001_),
    .X(_3004_));
 sky130_fd_sc_hd__nand2_1 _5975_ (.A(_3002_),
    .B(_3004_),
    .Y(_3005_));
 sky130_fd_sc_hd__or2_1 _5976_ (.A(_3000_),
    .B(_3005_),
    .X(_3006_));
 sky130_fd_sc_hd__a21oi_1 _5977_ (.A1(_3000_),
    .A2(_3005_),
    .B1(net2337),
    .Y(_3007_));
 sky130_fd_sc_hd__a32o_1 _5978_ (.A1(net204),
    .A2(_2732_),
    .A3(_2756_),
    .B1(_2986_),
    .B2(_2727_),
    .X(_3008_));
 sky130_fd_sc_hd__a221o_1 _5979_ (.A1(_1771_),
    .A2(_2769_),
    .B1(net350),
    .B2(_1768_),
    .C1(net211),
    .X(_3009_));
 sky130_fd_sc_hd__a22o_1 _5980_ (.A1(_1773_),
    .A2(net352),
    .B1(_3008_),
    .B2(net181),
    .X(_3010_));
 sky130_fd_sc_hd__mux4_1 _5981_ (.A0(_1708_),
    .A1(_1742_),
    .A2(_1770_),
    .A3(_1731_),
    .S0(_1681_),
    .S1(net189),
    .X(_3011_));
 sky130_fd_sc_hd__mux2_1 _5982_ (.A0(_2911_),
    .A1(_3011_),
    .S(net199),
    .X(_3012_));
 sky130_fd_sc_hd__o21ai_1 _5983_ (.A1(net197),
    .A2(_1846_),
    .B1(net202),
    .Y(_3013_));
 sky130_fd_sc_hd__o211ai_1 _5984_ (.A1(net202),
    .A2(_3012_),
    .B1(_3013_),
    .C1(_2775_),
    .Y(_3014_));
 sky130_fd_sc_hd__mux2_1 _5985_ (.A0(_2741_),
    .A1(_2749_),
    .S(net202),
    .X(_3015_));
 sky130_fd_sc_hd__a21bo_1 _5986_ (.A1(_2732_),
    .A2(_3015_),
    .B1_N(_3014_),
    .X(_3016_));
 sky130_fd_sc_hd__a22o_1 _5987_ (.A1(_3006_),
    .A2(_3007_),
    .B1(_3016_),
    .B2(net184),
    .X(_3017_));
 sky130_fd_sc_hd__a21oi_1 _5988_ (.A1(net2345),
    .A2(net211),
    .B1(net467),
    .Y(_3018_));
 sky130_fd_sc_hd__o31a_1 _5989_ (.A1(_3009_),
    .A2(_3010_),
    .A3(_3017_),
    .B1(_3018_),
    .X(_0852_));
 sky130_fd_sc_hd__xnor2_1 _5990_ (.A(_1792_),
    .B(net354),
    .Y(_3019_));
 sky130_fd_sc_hd__and2_1 _5991_ (.A(_1789_),
    .B(_3019_),
    .X(_3020_));
 sky130_fd_sc_hd__nand2_1 _5992_ (.A(_1789_),
    .B(_3019_),
    .Y(_3021_));
 sky130_fd_sc_hd__nor2_1 _5993_ (.A(_1789_),
    .B(_3019_),
    .Y(_3022_));
 sky130_fd_sc_hd__nor2_1 _5994_ (.A(_3020_),
    .B(_3022_),
    .Y(_3023_));
 sky130_fd_sc_hd__a21o_1 _5995_ (.A1(_3000_),
    .A2(_3002_),
    .B1(_3003_),
    .X(_3024_));
 sky130_fd_sc_hd__xor2_1 _5996_ (.A(_3023_),
    .B(_3024_),
    .X(_3025_));
 sky130_fd_sc_hd__mux4_1 _5997_ (.A0(_1708_),
    .A1(_1731_),
    .A2(_1770_),
    .A3(_1789_),
    .S0(net193),
    .S1(net188),
    .X(_3026_));
 sky130_fd_sc_hd__mux2_1 _5998_ (.A0(_2938_),
    .A1(_3026_),
    .S(net199),
    .X(_3027_));
 sky130_fd_sc_hd__nor2_1 _5999_ (.A(net201),
    .B(_3027_),
    .Y(_3028_));
 sky130_fd_sc_hd__a211o_1 _6000_ (.A1(net201),
    .A2(_2810_),
    .B1(_3028_),
    .C1(_2776_),
    .X(_3029_));
 sky130_fd_sc_hd__mux2_1 _6001_ (.A0(_2784_),
    .A1(_2821_),
    .S(net206),
    .X(_3030_));
 sky130_fd_sc_hd__a21bo_1 _6002_ (.A1(_2732_),
    .A2(_3030_),
    .B1_N(_3029_),
    .X(_3031_));
 sky130_fd_sc_hd__a221o_1 _6003_ (.A1(_1794_),
    .A2(net300),
    .B1(net350),
    .B2(_1792_),
    .C1(net211),
    .X(_3032_));
 sky130_fd_sc_hd__a22o_1 _6004_ (.A1(net352),
    .A2(_3023_),
    .B1(_3031_),
    .B2(net184),
    .X(_3033_));
 sky130_fd_sc_hd__nor2_1 _6005_ (.A(_3032_),
    .B(_3033_),
    .Y(_3034_));
 sky130_fd_sc_hd__a21oi_1 _6006_ (.A1(net204),
    .A2(_2791_),
    .B1(_2986_),
    .Y(_3035_));
 sky130_fd_sc_hd__nor2_2 _6007_ (.A(net203),
    .B(_2730_),
    .Y(_3036_));
 sky130_fd_sc_hd__nand2_1 _6008_ (.A(net204),
    .B(_2729_),
    .Y(_3037_));
 sky130_fd_sc_hd__o22a_1 _6009_ (.A1(_2728_),
    .A2(_3035_),
    .B1(_3037_),
    .B2(_2795_),
    .X(_3038_));
 sky130_fd_sc_hd__o22a_1 _6010_ (.A1(net302),
    .A2(_3025_),
    .B1(_3038_),
    .B2(net184),
    .X(_3039_));
 sky130_fd_sc_hd__a221oi_1 _6011_ (.A1(net2357),
    .A2(net211),
    .B1(_3034_),
    .B2(_3039_),
    .C1(net467),
    .Y(_0853_));
 sky130_fd_sc_hd__a21o_1 _6012_ (.A1(_3021_),
    .A2(_3024_),
    .B1(_3022_),
    .X(_3040_));
 sky130_fd_sc_hd__xnor2_1 _6013_ (.A(_1757_),
    .B(net354),
    .Y(_3041_));
 sky130_fd_sc_hd__nand2_1 _6014_ (.A(_1754_),
    .B(_3041_),
    .Y(_3042_));
 sky130_fd_sc_hd__nor2_1 _6015_ (.A(_1754_),
    .B(_3041_),
    .Y(_3043_));
 sky130_fd_sc_hd__or2_1 _6016_ (.A(_1754_),
    .B(_3041_),
    .X(_3044_));
 sky130_fd_sc_hd__nand2_1 _6017_ (.A(_3042_),
    .B(_3044_),
    .Y(_3045_));
 sky130_fd_sc_hd__xnor2_1 _6018_ (.A(_3040_),
    .B(_3045_),
    .Y(_3046_));
 sky130_fd_sc_hd__a21o_1 _6019_ (.A1(net204),
    .A2(_2849_),
    .B1(_2986_),
    .X(_3047_));
 sky130_fd_sc_hd__a22o_1 _6020_ (.A1(_2841_),
    .A2(_3036_),
    .B1(_3047_),
    .B2(_2727_),
    .X(_3048_));
 sky130_fd_sc_hd__a22o_1 _6021_ (.A1(_1758_),
    .A2(net300),
    .B1(net350),
    .B2(_1757_),
    .X(_3049_));
 sky130_fd_sc_hd__a22o_1 _6022_ (.A1(_1760_),
    .A2(net352),
    .B1(_3048_),
    .B2(net181),
    .X(_3050_));
 sky130_fd_sc_hd__nor3_1 _6023_ (.A(net210),
    .B(_3049_),
    .C(_3050_),
    .Y(_3051_));
 sky130_fd_sc_hd__mux4_1 _6024_ (.A0(_1731_),
    .A1(_1770_),
    .A2(_1789_),
    .A3(_1754_),
    .S0(net193),
    .S1(net189),
    .X(_3052_));
 sky130_fd_sc_hd__mux2_1 _6025_ (.A0(_2966_),
    .A1(_3052_),
    .S(net199),
    .X(_3053_));
 sky130_fd_sc_hd__or2_1 _6026_ (.A(net202),
    .B(_3053_),
    .X(_3054_));
 sky130_fd_sc_hd__o21ai_1 _6027_ (.A1(net207),
    .A2(_2828_),
    .B1(_3054_),
    .Y(_3055_));
 sky130_fd_sc_hd__mux2_1 _6028_ (.A0(_2835_),
    .A1(_2845_),
    .S(net202),
    .X(_3056_));
 sky130_fd_sc_hd__o2bb2a_1 _6029_ (.A1_N(_2732_),
    .A2_N(_3056_),
    .B1(_3055_),
    .B2(_2776_),
    .X(_3057_));
 sky130_fd_sc_hd__o22a_1 _6030_ (.A1(net2337),
    .A2(_3046_),
    .B1(_3057_),
    .B2(net181),
    .X(_3058_));
 sky130_fd_sc_hd__a221oi_1 _6031_ (.A1(_1759_),
    .A2(net210),
    .B1(_3051_),
    .B2(net2338),
    .C1(net467),
    .Y(_0854_));
 sky130_fd_sc_hd__xnor2_1 _6032_ (.A(_1781_),
    .B(net354),
    .Y(_3059_));
 sky130_fd_sc_hd__and2_1 _6033_ (.A(_1778_),
    .B(_3059_),
    .X(_3060_));
 sky130_fd_sc_hd__nand2_1 _6034_ (.A(_1778_),
    .B(_3059_),
    .Y(_3061_));
 sky130_fd_sc_hd__nor2_1 _6035_ (.A(_1778_),
    .B(_3059_),
    .Y(_3062_));
 sky130_fd_sc_hd__nor2_1 _6036_ (.A(_3060_),
    .B(_3062_),
    .Y(_3063_));
 sky130_fd_sc_hd__a21o_1 _6037_ (.A1(_3040_),
    .A2(_3042_),
    .B1(_3043_),
    .X(_3064_));
 sky130_fd_sc_hd__xor2_1 _6038_ (.A(_3063_),
    .B(_3064_),
    .X(_3065_));
 sky130_fd_sc_hd__mux4_1 _6039_ (.A0(_1754_),
    .A1(_1770_),
    .A2(_1778_),
    .A3(_1789_),
    .S0(net185),
    .S1(net192),
    .X(_3066_));
 sky130_fd_sc_hd__mux2_1 _6040_ (.A0(_2992_),
    .A1(_3066_),
    .S(net199),
    .X(_3067_));
 sky130_fd_sc_hd__a21o_1 _6041_ (.A1(net199),
    .A2(_2887_),
    .B1(net206),
    .X(_3068_));
 sky130_fd_sc_hd__o211ai_1 _6042_ (.A1(net201),
    .A2(_3067_),
    .B1(_3068_),
    .C1(_2775_),
    .Y(_3069_));
 sky130_fd_sc_hd__mux2_1 _6043_ (.A0(_2867_),
    .A1(_2896_),
    .S(net206),
    .X(_3070_));
 sky130_fd_sc_hd__a21bo_1 _6044_ (.A1(_2732_),
    .A2(_3070_),
    .B1_N(_3069_),
    .X(_3071_));
 sky130_fd_sc_hd__a221o_1 _6045_ (.A1(_1782_),
    .A2(net300),
    .B1(net350),
    .B2(_1781_),
    .C1(net210),
    .X(_3072_));
 sky130_fd_sc_hd__a22o_1 _6046_ (.A1(net352),
    .A2(_3063_),
    .B1(_3071_),
    .B2(net184),
    .X(_3073_));
 sky130_fd_sc_hd__a21oi_1 _6047_ (.A1(net204),
    .A2(_2871_),
    .B1(_2986_),
    .Y(_3074_));
 sky130_fd_sc_hd__o22a_1 _6048_ (.A1(_2874_),
    .A2(_3037_),
    .B1(_3074_),
    .B2(_2728_),
    .X(_3075_));
 sky130_fd_sc_hd__o22ai_1 _6049_ (.A1(net302),
    .A2(_3065_),
    .B1(_3075_),
    .B2(net184),
    .Y(_3076_));
 sky130_fd_sc_hd__a21oi_1 _6050_ (.A1(net2398),
    .A2(net210),
    .B1(net466),
    .Y(_3077_));
 sky130_fd_sc_hd__o31a_1 _6051_ (.A1(_3072_),
    .A2(_3073_),
    .A3(_3076_),
    .B1(_3077_),
    .X(_0855_));
 sky130_fd_sc_hd__a21o_1 _6052_ (.A1(_3061_),
    .A2(_3064_),
    .B1(_3062_),
    .X(_3078_));
 sky130_fd_sc_hd__xnor2_1 _6053_ (.A(_1812_),
    .B(net354),
    .Y(_3079_));
 sky130_fd_sc_hd__nand2_1 _6054_ (.A(_1815_),
    .B(_3079_),
    .Y(_3080_));
 sky130_fd_sc_hd__nor2_1 _6055_ (.A(_1815_),
    .B(_3079_),
    .Y(_3081_));
 sky130_fd_sc_hd__or2_1 _6056_ (.A(_1815_),
    .B(_3079_),
    .X(_3082_));
 sky130_fd_sc_hd__nand2_1 _6057_ (.A(_3080_),
    .B(_3082_),
    .Y(_3083_));
 sky130_fd_sc_hd__xnor2_1 _6058_ (.A(_3078_),
    .B(_3083_),
    .Y(_3084_));
 sky130_fd_sc_hd__a21oi_1 _6059_ (.A1(net204),
    .A2(_2909_),
    .B1(_2986_),
    .Y(_3085_));
 sky130_fd_sc_hd__a2bb2o_1 _6060_ (.A1_N(_2728_),
    .A2_N(_3085_),
    .B1(_3036_),
    .B2(_2908_),
    .X(_3086_));
 sky130_fd_sc_hd__a22o_1 _6061_ (.A1(_1816_),
    .A2(net300),
    .B1(net350),
    .B2(_1812_),
    .X(_3087_));
 sky130_fd_sc_hd__a22o_1 _6062_ (.A1(_1818_),
    .A2(net352),
    .B1(_3086_),
    .B2(net181),
    .X(_3088_));
 sky130_fd_sc_hd__nor3_1 _6063_ (.A(net210),
    .B(_3087_),
    .C(_3088_),
    .Y(_3089_));
 sky130_fd_sc_hd__mux4_1 _6064_ (.A0(_1754_),
    .A1(_1789_),
    .A2(_1815_),
    .A3(_1778_),
    .S0(net191),
    .S1(net188),
    .X(_3090_));
 sky130_fd_sc_hd__mux2_1 _6065_ (.A0(_3011_),
    .A1(_3090_),
    .S(net199),
    .X(_3091_));
 sky130_fd_sc_hd__or2_1 _6066_ (.A(net201),
    .B(_3091_),
    .X(_3092_));
 sky130_fd_sc_hd__o211a_1 _6067_ (.A1(net207),
    .A2(_2912_),
    .B1(_3092_),
    .C1(_2775_),
    .X(_3093_));
 sky130_fd_sc_hd__mux2_1 _6068_ (.A0(_2907_),
    .A1(_2914_),
    .S(net207),
    .X(_3094_));
 sky130_fd_sc_hd__a21oi_1 _6069_ (.A1(_2732_),
    .A2(_3094_),
    .B1(_3093_),
    .Y(_3095_));
 sky130_fd_sc_hd__o22a_1 _6070_ (.A1(net302),
    .A2(_3084_),
    .B1(_3095_),
    .B2(net181),
    .X(_3096_));
 sky130_fd_sc_hd__a221oi_1 _6071_ (.A1(_1817_),
    .A2(net210),
    .B1(_3089_),
    .B2(_3096_),
    .C1(net466),
    .Y(_0856_));
 sky130_fd_sc_hd__xnor2_1 _6072_ (.A(_1837_),
    .B(net354),
    .Y(_3097_));
 sky130_fd_sc_hd__and2_1 _6073_ (.A(_1834_),
    .B(_3097_),
    .X(_3098_));
 sky130_fd_sc_hd__nand2_1 _6074_ (.A(_1834_),
    .B(_3097_),
    .Y(_3099_));
 sky130_fd_sc_hd__nor2_1 _6075_ (.A(_1834_),
    .B(_3097_),
    .Y(_3100_));
 sky130_fd_sc_hd__nor2_1 _6076_ (.A(_3098_),
    .B(_3100_),
    .Y(_3101_));
 sky130_fd_sc_hd__a21o_1 _6077_ (.A1(_3078_),
    .A2(_3080_),
    .B1(_3081_),
    .X(_3102_));
 sky130_fd_sc_hd__xor2_1 _6078_ (.A(_3101_),
    .B(_3102_),
    .X(_3103_));
 sky130_fd_sc_hd__mux4_1 _6079_ (.A0(_1754_),
    .A1(_1778_),
    .A2(_1815_),
    .A3(_1834_),
    .S0(net192),
    .S1(net188),
    .X(_3104_));
 sky130_fd_sc_hd__or2_1 _6080_ (.A(net199),
    .B(_3026_),
    .X(_3105_));
 sky130_fd_sc_hd__o21ai_1 _6081_ (.A1(net196),
    .A2(_3104_),
    .B1(_3105_),
    .Y(_3106_));
 sky130_fd_sc_hd__mux2_1 _6082_ (.A0(_2940_),
    .A1(_3106_),
    .S(net206),
    .X(_3107_));
 sky130_fd_sc_hd__or2_1 _6083_ (.A(_2776_),
    .B(_3107_),
    .X(_3108_));
 sky130_fd_sc_hd__mux2_1 _6084_ (.A0(_2929_),
    .A1(_2942_),
    .S(net206),
    .X(_3109_));
 sky130_fd_sc_hd__a21bo_1 _6085_ (.A1(_2732_),
    .A2(_3109_),
    .B1_N(_3108_),
    .X(_3110_));
 sky130_fd_sc_hd__a221o_1 _6086_ (.A1(_1839_),
    .A2(net300),
    .B1(_2770_),
    .B2(_1837_),
    .C1(net210),
    .X(_3111_));
 sky130_fd_sc_hd__a22o_1 _6087_ (.A1(net352),
    .A2(_3101_),
    .B1(_3110_),
    .B2(net184),
    .X(_3112_));
 sky130_fd_sc_hd__o21a_1 _6088_ (.A1(net203),
    .A2(_2934_),
    .B1(_2987_),
    .X(_3113_));
 sky130_fd_sc_hd__a2bb2o_1 _6089_ (.A1_N(_2728_),
    .A2_N(_3113_),
    .B1(_3036_),
    .B2(_2931_),
    .X(_3114_));
 sky130_fd_sc_hd__a2bb2o_1 _6090_ (.A1_N(net302),
    .A2_N(_3103_),
    .B1(_3114_),
    .B2(net181),
    .X(_3115_));
 sky130_fd_sc_hd__a21oi_1 _6091_ (.A1(_1840_),
    .A2(net210),
    .B1(net466),
    .Y(_3116_));
 sky130_fd_sc_hd__o31a_1 _6092_ (.A1(_3111_),
    .A2(_3112_),
    .A3(_3115_),
    .B1(_3116_),
    .X(_0857_));
 sky130_fd_sc_hd__a21o_1 _6093_ (.A1(_3099_),
    .A2(_3102_),
    .B1(_3100_),
    .X(_3117_));
 sky130_fd_sc_hd__xnor2_1 _6094_ (.A(_1805_),
    .B(net354),
    .Y(_3118_));
 sky130_fd_sc_hd__nand2_1 _6095_ (.A(_1802_),
    .B(_3118_),
    .Y(_3119_));
 sky130_fd_sc_hd__or2_1 _6096_ (.A(_1802_),
    .B(_3118_),
    .X(_3120_));
 sky130_fd_sc_hd__nand2_1 _6097_ (.A(_3119_),
    .B(_3120_),
    .Y(_3121_));
 sky130_fd_sc_hd__xnor2_1 _6098_ (.A(_3117_),
    .B(_3121_),
    .Y(_3122_));
 sky130_fd_sc_hd__mux4_2 _6099_ (.A0(_1778_),
    .A1(_1815_),
    .A2(_1834_),
    .A3(_1802_),
    .S0(net192),
    .S1(net188),
    .X(_3123_));
 sky130_fd_sc_hd__mux2_1 _6100_ (.A0(_3052_),
    .A1(_3123_),
    .S(net200),
    .X(_3124_));
 sky130_fd_sc_hd__mux2_1 _6101_ (.A0(_2967_),
    .A1(_3124_),
    .S(net206),
    .X(_3125_));
 sky130_fd_sc_hd__mux2_1 _6102_ (.A0(_2956_),
    .A1(_2970_),
    .S(net207),
    .X(_3126_));
 sky130_fd_sc_hd__a22o_1 _6103_ (.A1(_2775_),
    .A2(_3125_),
    .B1(_3126_),
    .B2(_2732_),
    .X(_3127_));
 sky130_fd_sc_hd__o21a_1 _6104_ (.A1(_1802_),
    .A2(_1805_),
    .B1(net300),
    .X(_3128_));
 sky130_fd_sc_hd__a22o_1 _6105_ (.A1(_1806_),
    .A2(net352),
    .B1(_3127_),
    .B2(net184),
    .X(_3129_));
 sky130_fd_sc_hd__a2111o_1 _6106_ (.A1(_1805_),
    .A2(_2770_),
    .B1(net210),
    .C1(_3128_),
    .D1(_3129_),
    .X(_3130_));
 sky130_fd_sc_hd__a21oi_1 _6107_ (.A1(net204),
    .A2(_2960_),
    .B1(_2986_),
    .Y(_3131_));
 sky130_fd_sc_hd__o32a_1 _6108_ (.A1(net194),
    .A2(_2840_),
    .A3(_3037_),
    .B1(_3131_),
    .B2(_2728_),
    .X(_3132_));
 sky130_fd_sc_hd__o22ai_1 _6109_ (.A1(net302),
    .A2(_3122_),
    .B1(_3132_),
    .B2(net184),
    .Y(_3133_));
 sky130_fd_sc_hd__a21bo_1 _6110_ (.A1(net2373),
    .A2(_1805_),
    .B1_N(net210),
    .X(_3134_));
 sky130_fd_sc_hd__o211a_1 _6111_ (.A1(_3130_),
    .A2(_3133_),
    .B1(net2374),
    .C1(net446),
    .X(_0858_));
 sky130_fd_sc_hd__xnor2_1 _6112_ (.A(_1826_),
    .B(net353),
    .Y(_3135_));
 sky130_fd_sc_hd__and2_1 _6113_ (.A(_1823_),
    .B(_3135_),
    .X(_3136_));
 sky130_fd_sc_hd__nand2_1 _6114_ (.A(_1823_),
    .B(_3135_),
    .Y(_3137_));
 sky130_fd_sc_hd__nor2_1 _6115_ (.A(_1823_),
    .B(_3135_),
    .Y(_3138_));
 sky130_fd_sc_hd__nor2_1 _6116_ (.A(_3136_),
    .B(_3138_),
    .Y(_3139_));
 sky130_fd_sc_hd__a21bo_1 _6117_ (.A1(_3117_),
    .A2(_3119_),
    .B1_N(_3120_),
    .X(_3140_));
 sky130_fd_sc_hd__nand2_1 _6118_ (.A(_3139_),
    .B(_3140_),
    .Y(_3141_));
 sky130_fd_sc_hd__or2_1 _6119_ (.A(_3139_),
    .B(_3140_),
    .X(_3142_));
 sky130_fd_sc_hd__a21oi_1 _6120_ (.A1(_3141_),
    .A2(_3142_),
    .B1(net301),
    .Y(_3143_));
 sky130_fd_sc_hd__mux4_1 _6121_ (.A0(_1802_),
    .A1(_1815_),
    .A2(_1823_),
    .A3(_1834_),
    .S0(net185),
    .S1(net192),
    .X(_3144_));
 sky130_fd_sc_hd__mux2_1 _6122_ (.A0(_3066_),
    .A1(_3144_),
    .S(net198),
    .X(_3145_));
 sky130_fd_sc_hd__mux2_1 _6123_ (.A0(_2993_),
    .A1(_3145_),
    .S(net205),
    .X(_3146_));
 sky130_fd_sc_hd__a221o_1 _6124_ (.A1(_1827_),
    .A2(net299),
    .B1(net349),
    .B2(_1826_),
    .C1(net209),
    .X(_3147_));
 sky130_fd_sc_hd__a221o_1 _6125_ (.A1(net351),
    .A2(_3139_),
    .B1(_3146_),
    .B2(_2777_),
    .C1(_3147_),
    .X(_3148_));
 sky130_fd_sc_hd__nor2_2 _6126_ (.A(_1594_),
    .B(net183),
    .Y(_3149_));
 sky130_fd_sc_hd__nor2_4 _6127_ (.A(_2728_),
    .B(_3149_),
    .Y(_3150_));
 sky130_fd_sc_hd__or2_2 _6128_ (.A(_2728_),
    .B(_3149_),
    .X(_3151_));
 sky130_fd_sc_hd__nor2_2 _6129_ (.A(net180),
    .B(_2730_),
    .Y(_3152_));
 sky130_fd_sc_hd__or2_1 _6130_ (.A(_3150_),
    .B(_3152_),
    .X(_3153_));
 sky130_fd_sc_hd__a21o_1 _6131_ (.A1(_2983_),
    .A2(_3036_),
    .B1(_3153_),
    .X(_3154_));
 sky130_fd_sc_hd__mux2_1 _6132_ (.A0(_2981_),
    .A1(_2995_),
    .S(net205),
    .X(_3155_));
 sky130_fd_sc_hd__o21a_1 _6133_ (.A1(net180),
    .A2(_3155_),
    .B1(_3154_),
    .X(_3156_));
 sky130_fd_sc_hd__a21oi_1 _6134_ (.A1(_1828_),
    .A2(net209),
    .B1(net461),
    .Y(_3157_));
 sky130_fd_sc_hd__o31a_1 _6135_ (.A1(_3143_),
    .A2(_3148_),
    .A3(_3156_),
    .B1(_3157_),
    .X(_0859_));
 sky130_fd_sc_hd__a21o_1 _6136_ (.A1(_3137_),
    .A2(_3140_),
    .B1(_3138_),
    .X(_3158_));
 sky130_fd_sc_hd__xnor2_1 _6137_ (.A(_1511_),
    .B(net353),
    .Y(_3159_));
 sky130_fd_sc_hd__nand2_1 _6138_ (.A(_1513_),
    .B(_3159_),
    .Y(_3160_));
 sky130_fd_sc_hd__nor2_1 _6139_ (.A(_1513_),
    .B(_3159_),
    .Y(_3161_));
 sky130_fd_sc_hd__or2_1 _6140_ (.A(_1513_),
    .B(_3159_),
    .X(_3162_));
 sky130_fd_sc_hd__nand2_1 _6141_ (.A(_3160_),
    .B(_3162_),
    .Y(_3163_));
 sky130_fd_sc_hd__xnor2_1 _6142_ (.A(_3158_),
    .B(_3163_),
    .Y(_3164_));
 sky130_fd_sc_hd__mux4_1 _6143_ (.A0(_1513_),
    .A1(_1802_),
    .A2(_1823_),
    .A3(_1834_),
    .S0(net185),
    .S1(net190),
    .X(_3165_));
 sky130_fd_sc_hd__mux2_1 _6144_ (.A0(_3090_),
    .A1(_3165_),
    .S(net199),
    .X(_3166_));
 sky130_fd_sc_hd__mux2_1 _6145_ (.A0(_3012_),
    .A1(_3166_),
    .S(net206),
    .X(_3167_));
 sky130_fd_sc_hd__a31o_1 _6146_ (.A1(net206),
    .A2(net199),
    .A3(_1847_),
    .B1(net184),
    .X(_3168_));
 sky130_fd_sc_hd__o211a_1 _6147_ (.A1(net181),
    .A2(_3167_),
    .B1(_3168_),
    .C1(_2775_),
    .X(_3169_));
 sky130_fd_sc_hd__a221o_1 _6148_ (.A1(_1514_),
    .A2(net299),
    .B1(net349),
    .B2(_1511_),
    .C1(net209),
    .X(_3170_));
 sky130_fd_sc_hd__a221o_1 _6149_ (.A1(_1516_),
    .A2(net351),
    .B1(_3152_),
    .B2(_2757_),
    .C1(_3170_),
    .X(_3171_));
 sky130_fd_sc_hd__o21ai_1 _6150_ (.A1(net180),
    .A2(_2757_),
    .B1(_3150_),
    .Y(_3172_));
 sky130_fd_sc_hd__o21ai_1 _6151_ (.A1(net301),
    .A2(_3164_),
    .B1(_3172_),
    .Y(_3173_));
 sky130_fd_sc_hd__a21oi_1 _6152_ (.A1(_1515_),
    .A2(net209),
    .B1(net461),
    .Y(_3174_));
 sky130_fd_sc_hd__o31a_1 _6153_ (.A1(_3169_),
    .A2(_3171_),
    .A3(_3173_),
    .B1(_3174_),
    .X(_0860_));
 sky130_fd_sc_hd__xnor2_2 _6154_ (.A(_1526_),
    .B(net353),
    .Y(_3175_));
 sky130_fd_sc_hd__nand2_1 _6155_ (.A(_1521_),
    .B(_3175_),
    .Y(_3176_));
 sky130_fd_sc_hd__nor2_1 _6156_ (.A(_1521_),
    .B(_3175_),
    .Y(_3177_));
 sky130_fd_sc_hd__xor2_1 _6157_ (.A(_1521_),
    .B(_3175_),
    .X(_3178_));
 sky130_fd_sc_hd__a21o_1 _6158_ (.A1(_3158_),
    .A2(_3160_),
    .B1(_3161_),
    .X(_3179_));
 sky130_fd_sc_hd__xor2_1 _6159_ (.A(_3178_),
    .B(_3179_),
    .X(_3180_));
 sky130_fd_sc_hd__mux4_1 _6160_ (.A0(_1513_),
    .A1(_1521_),
    .A2(_1802_),
    .A3(_1823_),
    .S0(net192),
    .S1(net185),
    .X(_3181_));
 sky130_fd_sc_hd__mux2_1 _6161_ (.A0(_3104_),
    .A1(_3181_),
    .S(net198),
    .X(_3182_));
 sky130_fd_sc_hd__mux2_1 _6162_ (.A0(_3027_),
    .A1(_3182_),
    .S(net206),
    .X(_3183_));
 sky130_fd_sc_hd__nand2_1 _6163_ (.A(net181),
    .B(_2811_),
    .Y(_3184_));
 sky130_fd_sc_hd__o211a_1 _6164_ (.A1(net181),
    .A2(_3183_),
    .B1(_3184_),
    .C1(_2775_),
    .X(_3185_));
 sky130_fd_sc_hd__a221o_1 _6165_ (.A1(_1527_),
    .A2(net299),
    .B1(net349),
    .B2(_1526_),
    .C1(net209),
    .X(_3186_));
 sky130_fd_sc_hd__a221o_1 _6166_ (.A1(_2797_),
    .A2(_3152_),
    .B1(_3178_),
    .B2(net351),
    .C1(_3186_),
    .X(_3187_));
 sky130_fd_sc_hd__o21ai_1 _6167_ (.A1(net180),
    .A2(_2792_),
    .B1(_3150_),
    .Y(_3188_));
 sky130_fd_sc_hd__o21ai_1 _6168_ (.A1(net301),
    .A2(_3180_),
    .B1(_3188_),
    .Y(_3189_));
 sky130_fd_sc_hd__a21bo_1 _6169_ (.A1(_1521_),
    .A2(_1526_),
    .B1_N(net209),
    .X(_3190_));
 sky130_fd_sc_hd__o311a_1 _6170_ (.A1(_3185_),
    .A2(_3187_),
    .A3(_3189_),
    .B1(_3190_),
    .C1(net434),
    .X(_0861_));
 sky130_fd_sc_hd__a21o_1 _6171_ (.A1(_3176_),
    .A2(_3179_),
    .B1(_3177_),
    .X(_3191_));
 sky130_fd_sc_hd__xnor2_1 _6172_ (.A(_1536_),
    .B(net353),
    .Y(_3192_));
 sky130_fd_sc_hd__nand2_1 _6173_ (.A(_1533_),
    .B(_3192_),
    .Y(_3193_));
 sky130_fd_sc_hd__nor2_1 _6174_ (.A(_1533_),
    .B(_3192_),
    .Y(_3194_));
 sky130_fd_sc_hd__or2_1 _6175_ (.A(_1533_),
    .B(_3192_),
    .X(_3195_));
 sky130_fd_sc_hd__nand2_1 _6176_ (.A(_3193_),
    .B(_3195_),
    .Y(_3196_));
 sky130_fd_sc_hd__xnor2_1 _6177_ (.A(_3191_),
    .B(_3196_),
    .Y(_3197_));
 sky130_fd_sc_hd__mux4_1 _6178_ (.A0(_1513_),
    .A1(_1533_),
    .A2(_1823_),
    .A3(_1521_),
    .S0(net188),
    .S1(net190),
    .X(_3198_));
 sky130_fd_sc_hd__mux2_1 _6179_ (.A0(_3123_),
    .A1(_3198_),
    .S(net200),
    .X(_3199_));
 sky130_fd_sc_hd__mux2_1 _6180_ (.A0(_3053_),
    .A1(_3199_),
    .S(net205),
    .X(_3200_));
 sky130_fd_sc_hd__a21boi_1 _6181_ (.A1(_2775_),
    .A2(_3200_),
    .B1_N(_2847_),
    .Y(_3201_));
 sky130_fd_sc_hd__a22o_1 _6182_ (.A1(_1594_),
    .A2(_2727_),
    .B1(_2828_),
    .B2(_2829_),
    .X(_3202_));
 sky130_fd_sc_hd__a221o_1 _6183_ (.A1(_1538_),
    .A2(net299),
    .B1(net349),
    .B2(_1536_),
    .C1(net209),
    .X(_3203_));
 sky130_fd_sc_hd__a221o_1 _6184_ (.A1(_1540_),
    .A2(net351),
    .B1(_3202_),
    .B2(net180),
    .C1(_3203_),
    .X(_3204_));
 sky130_fd_sc_hd__o21ba_1 _6185_ (.A1(_2851_),
    .A2(_3149_),
    .B1_N(_3204_),
    .X(_3205_));
 sky130_fd_sc_hd__o221a_1 _6186_ (.A1(net301),
    .A2(_3197_),
    .B1(_3201_),
    .B2(net180),
    .C1(_3205_),
    .X(_3206_));
 sky130_fd_sc_hd__a211oi_1 _6187_ (.A1(_1537_),
    .A2(net209),
    .B1(_3206_),
    .C1(net462),
    .Y(_0862_));
 sky130_fd_sc_hd__xnor2_1 _6188_ (.A(_1548_),
    .B(net353),
    .Y(_3207_));
 sky130_fd_sc_hd__and2_1 _6189_ (.A(_1545_),
    .B(_3207_),
    .X(_3208_));
 sky130_fd_sc_hd__nand2_1 _6190_ (.A(_1545_),
    .B(_3207_),
    .Y(_3209_));
 sky130_fd_sc_hd__nor2_1 _6191_ (.A(_1545_),
    .B(_3207_),
    .Y(_3210_));
 sky130_fd_sc_hd__nor2_1 _6192_ (.A(_3208_),
    .B(_3210_),
    .Y(_3211_));
 sky130_fd_sc_hd__a21o_1 _6193_ (.A1(_3191_),
    .A2(_3193_),
    .B1(_3194_),
    .X(_3212_));
 sky130_fd_sc_hd__xor2_1 _6194_ (.A(_3211_),
    .B(_3212_),
    .X(_3213_));
 sky130_fd_sc_hd__mux4_1 _6195_ (.A0(_1513_),
    .A1(_1521_),
    .A2(_1533_),
    .A3(_1545_),
    .S0(net192),
    .S1(net188),
    .X(_3214_));
 sky130_fd_sc_hd__mux2_1 _6196_ (.A0(_3144_),
    .A1(_3214_),
    .S(net198),
    .X(_3215_));
 sky130_fd_sc_hd__mux2_1 _6197_ (.A0(_3067_),
    .A1(_3215_),
    .S(net206),
    .X(_3216_));
 sky130_fd_sc_hd__mux2_1 _6198_ (.A0(_2888_),
    .A1(_3216_),
    .S(net184),
    .X(_3217_));
 sky130_fd_sc_hd__a221o_1 _6199_ (.A1(_1549_),
    .A2(net299),
    .B1(net349),
    .B2(_1548_),
    .C1(net209),
    .X(_3218_));
 sky130_fd_sc_hd__a221o_1 _6200_ (.A1(_2876_),
    .A2(_3152_),
    .B1(_3211_),
    .B2(net351),
    .C1(_3218_),
    .X(_3219_));
 sky130_fd_sc_hd__o21ai_1 _6201_ (.A1(net180),
    .A2(_2872_),
    .B1(_3150_),
    .Y(_3220_));
 sky130_fd_sc_hd__a21oi_1 _6202_ (.A1(_2775_),
    .A2(_3217_),
    .B1(_3219_),
    .Y(_3221_));
 sky130_fd_sc_hd__o211a_1 _6203_ (.A1(net301),
    .A2(_3213_),
    .B1(_3220_),
    .C1(_3221_),
    .X(_3222_));
 sky130_fd_sc_hd__a211oi_1 _6204_ (.A1(net2367),
    .A2(net209),
    .B1(_3222_),
    .C1(net462),
    .Y(_0863_));
 sky130_fd_sc_hd__a21o_1 _6205_ (.A1(_3209_),
    .A2(_3212_),
    .B1(_3210_),
    .X(_3223_));
 sky130_fd_sc_hd__xnor2_1 _6206_ (.A(_1618_),
    .B(_2760_),
    .Y(_3224_));
 sky130_fd_sc_hd__nand2_1 _6207_ (.A(_1621_),
    .B(_3224_),
    .Y(_3225_));
 sky130_fd_sc_hd__nor2_1 _6208_ (.A(_1621_),
    .B(_3224_),
    .Y(_3226_));
 sky130_fd_sc_hd__or2_1 _6209_ (.A(_1621_),
    .B(_3224_),
    .X(_3227_));
 sky130_fd_sc_hd__nand2_1 _6210_ (.A(_3225_),
    .B(_3227_),
    .Y(_3228_));
 sky130_fd_sc_hd__xnor2_1 _6211_ (.A(_3223_),
    .B(_3228_),
    .Y(_3229_));
 sky130_fd_sc_hd__nor2_1 _6212_ (.A(net301),
    .B(_3229_),
    .Y(_3230_));
 sky130_fd_sc_hd__o32a_1 _6213_ (.A1(net204),
    .A2(_2908_),
    .A3(_3150_),
    .B1(_2910_),
    .B2(net182),
    .X(_3231_));
 sky130_fd_sc_hd__a21o_1 _6214_ (.A1(_2829_),
    .A2(_2912_),
    .B1(_2777_),
    .X(_3232_));
 sky130_fd_sc_hd__mux4_1 _6215_ (.A0(_1521_),
    .A1(_1533_),
    .A2(_1545_),
    .A3(_1621_),
    .S0(net192),
    .S1(net188),
    .X(_3233_));
 sky130_fd_sc_hd__mux2_1 _6216_ (.A0(_3165_),
    .A1(_3233_),
    .S(net198),
    .X(_3234_));
 sky130_fd_sc_hd__or3_1 _6217_ (.A(net201),
    .B(net180),
    .C(_3234_),
    .X(_3235_));
 sky130_fd_sc_hd__o211a_1 _6218_ (.A1(net206),
    .A2(_3091_),
    .B1(_3232_),
    .C1(_3235_),
    .X(_3236_));
 sky130_fd_sc_hd__a221o_1 _6219_ (.A1(_1622_),
    .A2(net299),
    .B1(net349),
    .B2(_1619_),
    .C1(net209),
    .X(_3237_));
 sky130_fd_sc_hd__a22o_1 _6220_ (.A1(_1624_),
    .A2(net351),
    .B1(_3153_),
    .B2(_3231_),
    .X(_3238_));
 sky130_fd_sc_hd__a21oi_1 _6221_ (.A1(_1623_),
    .A2(net209),
    .B1(net462),
    .Y(_3239_));
 sky130_fd_sc_hd__o41a_1 _6222_ (.A1(_3230_),
    .A2(_3236_),
    .A3(_3237_),
    .A4(_3238_),
    .B1(_3239_),
    .X(_0864_));
 sky130_fd_sc_hd__xnor2_1 _6223_ (.A(_1643_),
    .B(net353),
    .Y(_3240_));
 sky130_fd_sc_hd__and2_1 _6224_ (.A(_1640_),
    .B(_3240_),
    .X(_3241_));
 sky130_fd_sc_hd__nand2_1 _6225_ (.A(_1640_),
    .B(_3240_),
    .Y(_3242_));
 sky130_fd_sc_hd__nor2_1 _6226_ (.A(_1640_),
    .B(_3240_),
    .Y(_3243_));
 sky130_fd_sc_hd__nor2_1 _6227_ (.A(_3241_),
    .B(_3243_),
    .Y(_3244_));
 sky130_fd_sc_hd__a21o_1 _6228_ (.A1(_3223_),
    .A2(_3225_),
    .B1(_3226_),
    .X(_3245_));
 sky130_fd_sc_hd__xor2_1 _6229_ (.A(_3244_),
    .B(_3245_),
    .X(_3246_));
 sky130_fd_sc_hd__o21ai_1 _6230_ (.A1(net180),
    .A2(_2935_),
    .B1(_3150_),
    .Y(_3247_));
 sky130_fd_sc_hd__a221o_1 _6231_ (.A1(_1645_),
    .A2(net299),
    .B1(net349),
    .B2(_1643_),
    .C1(net209),
    .X(_3248_));
 sky130_fd_sc_hd__a21oi_1 _6232_ (.A1(net351),
    .A2(_3244_),
    .B1(_3248_),
    .Y(_3249_));
 sky130_fd_sc_hd__mux4_1 _6233_ (.A0(_1533_),
    .A1(_1545_),
    .A2(_1621_),
    .A3(_1640_),
    .S0(net192),
    .S1(net188),
    .X(_3250_));
 sky130_fd_sc_hd__mux2_1 _6234_ (.A0(_3181_),
    .A1(_3250_),
    .S(net198),
    .X(_3251_));
 sky130_fd_sc_hd__nand2_1 _6235_ (.A(net205),
    .B(_3251_),
    .Y(_3252_));
 sky130_fd_sc_hd__o211a_1 _6236_ (.A1(net205),
    .A2(_3106_),
    .B1(_3252_),
    .C1(net183),
    .X(_3253_));
 sky130_fd_sc_hd__o31a_1 _6237_ (.A1(net201),
    .A2(_2776_),
    .A3(_2940_),
    .B1(_2778_),
    .X(_3254_));
 sky130_fd_sc_hd__o22a_1 _6238_ (.A1(net301),
    .A2(_3246_),
    .B1(_3253_),
    .B2(_3254_),
    .X(_3255_));
 sky130_fd_sc_hd__o211a_1 _6239_ (.A1(net180),
    .A2(_2933_),
    .B1(_3249_),
    .C1(_3255_),
    .X(_3256_));
 sky130_fd_sc_hd__a221oi_2 _6240_ (.A1(_1646_),
    .A2(net209),
    .B1(_3247_),
    .B2(_3256_),
    .C1(net462),
    .Y(_0865_));
 sky130_fd_sc_hd__a21o_1 _6241_ (.A1(_3242_),
    .A2(_3245_),
    .B1(_3243_),
    .X(_3257_));
 sky130_fd_sc_hd__xnor2_1 _6242_ (.A(_1608_),
    .B(net353),
    .Y(_3258_));
 sky130_fd_sc_hd__nand2_1 _6243_ (.A(_1605_),
    .B(_3258_),
    .Y(_3259_));
 sky130_fd_sc_hd__nor2_1 _6244_ (.A(_1605_),
    .B(_3258_),
    .Y(_3260_));
 sky130_fd_sc_hd__inv_2 _6245_ (.A(_3260_),
    .Y(_3261_));
 sky130_fd_sc_hd__nand2_1 _6246_ (.A(_3259_),
    .B(_3261_),
    .Y(_3262_));
 sky130_fd_sc_hd__xnor2_1 _6247_ (.A(_3257_),
    .B(_3262_),
    .Y(_3263_));
 sky130_fd_sc_hd__mux4_1 _6248_ (.A0(_1545_),
    .A1(_1621_),
    .A2(_1640_),
    .A3(_1605_),
    .S0(_1680_),
    .S1(net189),
    .X(_3264_));
 sky130_fd_sc_hd__mux2_1 _6249_ (.A0(_3198_),
    .A1(_3264_),
    .S(net198),
    .X(_3265_));
 sky130_fd_sc_hd__mux2_1 _6250_ (.A0(_3124_),
    .A1(_3265_),
    .S(net207),
    .X(_3266_));
 sky130_fd_sc_hd__nor2_1 _6251_ (.A(net182),
    .B(_3266_),
    .Y(_3267_));
 sky130_fd_sc_hd__a211o_1 _6252_ (.A1(net182),
    .A2(_2968_),
    .B1(_3267_),
    .C1(_2776_),
    .X(_3268_));
 sky130_fd_sc_hd__a21oi_1 _6253_ (.A1(net183),
    .A2(_2961_),
    .B1(_3151_),
    .Y(_3269_));
 sky130_fd_sc_hd__a221o_1 _6254_ (.A1(_1609_),
    .A2(net299),
    .B1(net349),
    .B2(_1608_),
    .C1(net208),
    .X(_3270_));
 sky130_fd_sc_hd__a221o_1 _6255_ (.A1(_1611_),
    .A2(net351),
    .B1(_2959_),
    .B2(net183),
    .C1(_3270_),
    .X(_3271_));
 sky130_fd_sc_hd__o21ai_1 _6256_ (.A1(net301),
    .A2(_3263_),
    .B1(_3268_),
    .Y(_3272_));
 sky130_fd_sc_hd__a21oi_1 _6257_ (.A1(_1610_),
    .A2(net208),
    .B1(net462),
    .Y(_3273_));
 sky130_fd_sc_hd__o31a_1 _6258_ (.A1(_3269_),
    .A2(_3271_),
    .A3(_3272_),
    .B1(_3273_),
    .X(_0866_));
 sky130_fd_sc_hd__xnor2_1 _6259_ (.A(_1632_),
    .B(net353),
    .Y(_3274_));
 sky130_fd_sc_hd__and2_1 _6260_ (.A(_1629_),
    .B(_3274_),
    .X(_3275_));
 sky130_fd_sc_hd__nand2_1 _6261_ (.A(_1629_),
    .B(_3274_),
    .Y(_3276_));
 sky130_fd_sc_hd__nor2_1 _6262_ (.A(_1629_),
    .B(_3274_),
    .Y(_3277_));
 sky130_fd_sc_hd__nor2_1 _6263_ (.A(_3275_),
    .B(_3277_),
    .Y(_3278_));
 sky130_fd_sc_hd__a21o_1 _6264_ (.A1(_3257_),
    .A2(_3259_),
    .B1(_3260_),
    .X(_3279_));
 sky130_fd_sc_hd__nand2_1 _6265_ (.A(_3278_),
    .B(_3279_),
    .Y(_3280_));
 sky130_fd_sc_hd__or2_1 _6266_ (.A(_3278_),
    .B(_3279_),
    .X(_3281_));
 sky130_fd_sc_hd__a21oi_1 _6267_ (.A1(_3280_),
    .A2(_3281_),
    .B1(net301),
    .Y(_3282_));
 sky130_fd_sc_hd__mux4_1 _6268_ (.A0(_1605_),
    .A1(_1621_),
    .A2(_1629_),
    .A3(_1640_),
    .S0(net185),
    .S1(net192),
    .X(_3283_));
 sky130_fd_sc_hd__mux2_1 _6269_ (.A0(_3214_),
    .A1(_3283_),
    .S(net198),
    .X(_3284_));
 sky130_fd_sc_hd__or2_1 _6270_ (.A(net203),
    .B(_3284_),
    .X(_3285_));
 sky130_fd_sc_hd__o211a_1 _6271_ (.A1(net205),
    .A2(_3145_),
    .B1(_3285_),
    .C1(_2775_),
    .X(_3286_));
 sky130_fd_sc_hd__a221o_1 _6272_ (.A1(_1633_),
    .A2(net299),
    .B1(net349),
    .B2(_1632_),
    .C1(net208),
    .X(_3287_));
 sky130_fd_sc_hd__a221o_1 _6273_ (.A1(_1594_),
    .A2(_2727_),
    .B1(_2829_),
    .B2(_2993_),
    .C1(net183),
    .X(_3288_));
 sky130_fd_sc_hd__o31a_1 _6274_ (.A1(net180),
    .A2(_2985_),
    .A3(_3286_),
    .B1(_3288_),
    .X(_3289_));
 sky130_fd_sc_hd__a221o_1 _6275_ (.A1(_2988_),
    .A2(_3150_),
    .B1(_3278_),
    .B2(net351),
    .C1(_3287_),
    .X(_3290_));
 sky130_fd_sc_hd__a21oi_1 _6276_ (.A1(_1634_),
    .A2(net208),
    .B1(net462),
    .Y(_3291_));
 sky130_fd_sc_hd__o31a_1 _6277_ (.A1(_3282_),
    .A2(_3289_),
    .A3(_3290_),
    .B1(_3291_),
    .X(_0867_));
 sky130_fd_sc_hd__a21o_1 _6278_ (.A1(_3276_),
    .A2(_3279_),
    .B1(_3277_),
    .X(_3292_));
 sky130_fd_sc_hd__xnor2_1 _6279_ (.A(_1484_),
    .B(net353),
    .Y(_3293_));
 sky130_fd_sc_hd__nor2_1 _6280_ (.A(_1487_),
    .B(_3293_),
    .Y(_3294_));
 sky130_fd_sc_hd__nand2_1 _6281_ (.A(_1487_),
    .B(_3293_),
    .Y(_3295_));
 sky130_fd_sc_hd__and2b_1 _6282_ (.A_N(_3294_),
    .B(_3295_),
    .X(_3296_));
 sky130_fd_sc_hd__xor2_1 _6283_ (.A(_3292_),
    .B(_3296_),
    .X(_3297_));
 sky130_fd_sc_hd__mux4_1 _6284_ (.A0(_1487_),
    .A1(_1605_),
    .A2(_1629_),
    .A3(_1640_),
    .S0(net185),
    .S1(net190),
    .X(_3298_));
 sky130_fd_sc_hd__mux2_1 _6285_ (.A0(_3233_),
    .A1(_3298_),
    .S(net198),
    .X(_3299_));
 sky130_fd_sc_hd__mux2_1 _6286_ (.A0(_3166_),
    .A1(_3299_),
    .S(net206),
    .X(_3300_));
 sky130_fd_sc_hd__o2bb2a_1 _6287_ (.A1_N(_2778_),
    .A2_N(_3014_),
    .B1(_3300_),
    .B2(net182),
    .X(_3301_));
 sky130_fd_sc_hd__a221o_1 _6288_ (.A1(_1488_),
    .A2(net351),
    .B1(net349),
    .B2(_1484_),
    .C1(net299),
    .X(_3302_));
 sky130_fd_sc_hd__o21a_1 _6289_ (.A1(_1484_),
    .A2(_1487_),
    .B1(_3302_),
    .X(_3303_));
 sky130_fd_sc_hd__o211a_1 _6290_ (.A1(net203),
    .A2(net180),
    .B1(_2727_),
    .C1(_1594_),
    .X(_3304_));
 sky130_fd_sc_hd__a31o_1 _6291_ (.A1(net204),
    .A2(_2756_),
    .A3(_3153_),
    .B1(_3301_),
    .X(_3305_));
 sky130_fd_sc_hd__or4_1 _6292_ (.A(net208),
    .B(_3303_),
    .C(_3304_),
    .D(_3305_),
    .X(_3306_));
 sky130_fd_sc_hd__o21ba_1 _6293_ (.A1(net301),
    .A2(_3297_),
    .B1_N(_3306_),
    .X(_3307_));
 sky130_fd_sc_hd__a211oi_1 _6294_ (.A1(net2331),
    .A2(net208),
    .B1(_3307_),
    .C1(net462),
    .Y(_0868_));
 sky130_fd_sc_hd__xnor2_1 _6295_ (.A(_1462_),
    .B(net353),
    .Y(_3308_));
 sky130_fd_sc_hd__and2_1 _6296_ (.A(_1438_),
    .B(_3308_),
    .X(_3309_));
 sky130_fd_sc_hd__nand2_1 _6297_ (.A(_1438_),
    .B(_3308_),
    .Y(_3310_));
 sky130_fd_sc_hd__nor2_1 _6298_ (.A(_1438_),
    .B(_3308_),
    .Y(_3311_));
 sky130_fd_sc_hd__nor2_1 _6299_ (.A(_3309_),
    .B(_3311_),
    .Y(_3312_));
 sky130_fd_sc_hd__a21o_1 _6300_ (.A1(_3292_),
    .A2(_3295_),
    .B1(_3294_),
    .X(_3313_));
 sky130_fd_sc_hd__xor2_1 _6301_ (.A(_3312_),
    .B(_3313_),
    .X(_3314_));
 sky130_fd_sc_hd__nand2_1 _6302_ (.A(net201),
    .B(_3182_),
    .Y(_3315_));
 sky130_fd_sc_hd__mux4_1 _6303_ (.A0(_1438_),
    .A1(_1487_),
    .A2(_1629_),
    .A3(_1605_),
    .S0(net190),
    .S1(net185),
    .X(_3316_));
 sky130_fd_sc_hd__mux2_1 _6304_ (.A0(_3250_),
    .A1(_3316_),
    .S(net198),
    .X(_3317_));
 sky130_fd_sc_hd__nand2_1 _6305_ (.A(net205),
    .B(_3317_),
    .Y(_3318_));
 sky130_fd_sc_hd__a32o_1 _6306_ (.A1(net183),
    .A2(_3315_),
    .A3(_3318_),
    .B1(_2778_),
    .B2(_3029_),
    .X(_3319_));
 sky130_fd_sc_hd__nand2_1 _6307_ (.A(_1721_),
    .B(_3035_),
    .Y(_3320_));
 sky130_fd_sc_hd__a221o_1 _6308_ (.A1(_1464_),
    .A2(net299),
    .B1(net349),
    .B2(_1462_),
    .C1(net208),
    .X(_3321_));
 sky130_fd_sc_hd__nor2_2 _6309_ (.A(net180),
    .B(_3037_),
    .Y(_3322_));
 sky130_fd_sc_hd__a221o_1 _6310_ (.A1(net351),
    .A2(_3312_),
    .B1(_3322_),
    .B2(_2796_),
    .C1(_3321_),
    .X(_3323_));
 sky130_fd_sc_hd__a21oi_1 _6311_ (.A1(_3150_),
    .A2(_3320_),
    .B1(_3323_),
    .Y(_3324_));
 sky130_fd_sc_hd__o211a_1 _6312_ (.A1(net301),
    .A2(_3314_),
    .B1(_3319_),
    .C1(_3324_),
    .X(_3325_));
 sky130_fd_sc_hd__a211oi_2 _6313_ (.A1(_1465_),
    .A2(net208),
    .B1(_3325_),
    .C1(net462),
    .Y(_0869_));
 sky130_fd_sc_hd__a21o_1 _6314_ (.A1(_3310_),
    .A2(_3313_),
    .B1(_3311_),
    .X(_3326_));
 sky130_fd_sc_hd__xnor2_1 _6315_ (.A(_1474_),
    .B(net353),
    .Y(_3327_));
 sky130_fd_sc_hd__nand2_1 _6316_ (.A(_1471_),
    .B(_3327_),
    .Y(_3328_));
 sky130_fd_sc_hd__nor2_1 _6317_ (.A(_1471_),
    .B(_3327_),
    .Y(_3329_));
 sky130_fd_sc_hd__or2_1 _6318_ (.A(_1471_),
    .B(_3327_),
    .X(_3330_));
 sky130_fd_sc_hd__nand2_1 _6319_ (.A(_3328_),
    .B(_3330_),
    .Y(_3331_));
 sky130_fd_sc_hd__xnor2_1 _6320_ (.A(_3326_),
    .B(_3331_),
    .Y(_3332_));
 sky130_fd_sc_hd__o21a_1 _6321_ (.A1(_2776_),
    .A2(_3055_),
    .B1(_3151_),
    .X(_3333_));
 sky130_fd_sc_hd__mux4_1 _6322_ (.A0(_1438_),
    .A1(_1471_),
    .A2(_1629_),
    .A3(_1487_),
    .S0(net193),
    .S1(net186),
    .X(_3334_));
 sky130_fd_sc_hd__mux2_1 _6323_ (.A0(_3264_),
    .A1(_3334_),
    .S(net198),
    .X(_3335_));
 sky130_fd_sc_hd__mux2_1 _6324_ (.A0(_3199_),
    .A1(_3335_),
    .S(net205),
    .X(_3336_));
 sky130_fd_sc_hd__a22o_1 _6325_ (.A1(_2841_),
    .A2(_3036_),
    .B1(_3336_),
    .B2(_2775_),
    .X(_3337_));
 sky130_fd_sc_hd__a221o_1 _6326_ (.A1(_1476_),
    .A2(net299),
    .B1(net349),
    .B2(_1474_),
    .C1(net208),
    .X(_3338_));
 sky130_fd_sc_hd__a221o_1 _6327_ (.A1(_1477_),
    .A2(net351),
    .B1(_3047_),
    .B2(_3150_),
    .C1(_3338_),
    .X(_3339_));
 sky130_fd_sc_hd__a21oi_1 _6328_ (.A1(net183),
    .A2(_3337_),
    .B1(_3339_),
    .Y(_3340_));
 sky130_fd_sc_hd__o221a_1 _6329_ (.A1(net301),
    .A2(_3332_),
    .B1(_3333_),
    .B2(net183),
    .C1(_3340_),
    .X(_3341_));
 sky130_fd_sc_hd__a211oi_1 _6330_ (.A1(_1475_),
    .A2(net208),
    .B1(_3341_),
    .C1(net464),
    .Y(_0870_));
 sky130_fd_sc_hd__xnor2_1 _6331_ (.A(_1498_),
    .B(net353),
    .Y(_3342_));
 sky130_fd_sc_hd__and2_1 _6332_ (.A(_1494_),
    .B(_3342_),
    .X(_3343_));
 sky130_fd_sc_hd__nand2_1 _6333_ (.A(_1494_),
    .B(_3342_),
    .Y(_3344_));
 sky130_fd_sc_hd__nor2_1 _6334_ (.A(_1494_),
    .B(_3342_),
    .Y(_3345_));
 sky130_fd_sc_hd__nor2_1 _6335_ (.A(_3343_),
    .B(_3345_),
    .Y(_3346_));
 sky130_fd_sc_hd__a21o_1 _6336_ (.A1(_3326_),
    .A2(_3328_),
    .B1(_3329_),
    .X(_3347_));
 sky130_fd_sc_hd__nand2_1 _6337_ (.A(_3346_),
    .B(_3347_),
    .Y(_3348_));
 sky130_fd_sc_hd__or2_1 _6338_ (.A(_3346_),
    .B(_3347_),
    .X(_3349_));
 sky130_fd_sc_hd__a21oi_1 _6339_ (.A1(_3348_),
    .A2(_3349_),
    .B1(net301),
    .Y(_3350_));
 sky130_fd_sc_hd__mux4_1 _6340_ (.A0(_1438_),
    .A1(_1487_),
    .A2(_1494_),
    .A3(_1471_),
    .S0(net190),
    .S1(net188),
    .X(_3351_));
 sky130_fd_sc_hd__mux2_1 _6341_ (.A0(_3283_),
    .A1(_3351_),
    .S(net198),
    .X(_3352_));
 sky130_fd_sc_hd__mux2_1 _6342_ (.A0(_3215_),
    .A1(_3352_),
    .S(net206),
    .X(_3353_));
 sky130_fd_sc_hd__o2bb2a_1 _6343_ (.A1_N(_2778_),
    .A2_N(_3069_),
    .B1(_3353_),
    .B2(net180),
    .X(_3354_));
 sky130_fd_sc_hd__a21oi_1 _6344_ (.A1(net183),
    .A2(_3074_),
    .B1(_3151_),
    .Y(_3355_));
 sky130_fd_sc_hd__a221o_1 _6345_ (.A1(_1499_),
    .A2(net299),
    .B1(net349),
    .B2(_1498_),
    .C1(net208),
    .X(_3356_));
 sky130_fd_sc_hd__a221o_1 _6346_ (.A1(_2875_),
    .A2(_3322_),
    .B1(_3346_),
    .B2(net351),
    .C1(_3356_),
    .X(_3357_));
 sky130_fd_sc_hd__a21oi_1 _6347_ (.A1(_1500_),
    .A2(net208),
    .B1(net462),
    .Y(_3358_));
 sky130_fd_sc_hd__o41a_1 _6348_ (.A1(_3350_),
    .A2(_3354_),
    .A3(_3355_),
    .A4(_3357_),
    .B1(_3358_),
    .X(_0871_));
 sky130_fd_sc_hd__a21o_1 _6349_ (.A1(_3344_),
    .A2(_3347_),
    .B1(_3345_),
    .X(_3359_));
 sky130_fd_sc_hd__xnor2_1 _6350_ (.A(_1569_),
    .B(net353),
    .Y(_3360_));
 sky130_fd_sc_hd__nand2_1 _6351_ (.A(_1572_),
    .B(_3360_),
    .Y(_3361_));
 sky130_fd_sc_hd__nor2_1 _6352_ (.A(_1572_),
    .B(_3360_),
    .Y(_3362_));
 sky130_fd_sc_hd__inv_2 _6353_ (.A(_3362_),
    .Y(_3363_));
 sky130_fd_sc_hd__a21oi_1 _6354_ (.A1(_3361_),
    .A2(_3363_),
    .B1(_3359_),
    .Y(_3364_));
 sky130_fd_sc_hd__and3_1 _6355_ (.A(_3359_),
    .B(_3361_),
    .C(_3363_),
    .X(_3365_));
 sky130_fd_sc_hd__o21ba_1 _6356_ (.A1(_3364_),
    .A2(_3365_),
    .B1_N(net301),
    .X(_3366_));
 sky130_fd_sc_hd__mux4_1 _6357_ (.A0(_1438_),
    .A1(_1471_),
    .A2(_1494_),
    .A3(_1572_),
    .S0(net192),
    .S1(net189),
    .X(_3367_));
 sky130_fd_sc_hd__mux2_1 _6358_ (.A0(_3298_),
    .A1(_3367_),
    .S(net198),
    .X(_3368_));
 sky130_fd_sc_hd__mux2_1 _6359_ (.A0(_3234_),
    .A1(_3368_),
    .S(net205),
    .X(_3369_));
 sky130_fd_sc_hd__o22a_1 _6360_ (.A1(_2777_),
    .A2(_3093_),
    .B1(_3369_),
    .B2(net182),
    .X(_3370_));
 sky130_fd_sc_hd__nand2_1 _6361_ (.A(net183),
    .B(_3085_),
    .Y(_3371_));
 sky130_fd_sc_hd__and3_1 _6362_ (.A(net183),
    .B(_2908_),
    .C(_3036_),
    .X(_3372_));
 sky130_fd_sc_hd__a221o_1 _6363_ (.A1(_1573_),
    .A2(net299),
    .B1(net349),
    .B2(_1569_),
    .C1(_2772_),
    .X(_3373_));
 sky130_fd_sc_hd__a221o_1 _6364_ (.A1(_1575_),
    .A2(net351),
    .B1(_3150_),
    .B2(_3371_),
    .C1(_3372_),
    .X(_3374_));
 sky130_fd_sc_hd__a21oi_1 _6365_ (.A1(_1574_),
    .A2(_2772_),
    .B1(net464),
    .Y(_3375_));
 sky130_fd_sc_hd__o41a_1 _6366_ (.A1(_3366_),
    .A2(_3370_),
    .A3(_3373_),
    .A4(_3374_),
    .B1(_3375_),
    .X(_0872_));
 sky130_fd_sc_hd__xnor2_1 _6367_ (.A(_1584_),
    .B(net353),
    .Y(_3376_));
 sky130_fd_sc_hd__nand2_1 _6368_ (.A(_1580_),
    .B(_3376_),
    .Y(_3377_));
 sky130_fd_sc_hd__nor2_1 _6369_ (.A(_1580_),
    .B(_3376_),
    .Y(_3378_));
 sky130_fd_sc_hd__or2_1 _6370_ (.A(_1580_),
    .B(_3376_),
    .X(_3379_));
 sky130_fd_sc_hd__nand2_1 _6371_ (.A(_3377_),
    .B(_3379_),
    .Y(_3380_));
 sky130_fd_sc_hd__a21o_1 _6372_ (.A1(_3359_),
    .A2(_3361_),
    .B1(_3362_),
    .X(_3381_));
 sky130_fd_sc_hd__xnor2_1 _6373_ (.A(_3380_),
    .B(_3381_),
    .Y(_3382_));
 sky130_fd_sc_hd__mux4_1 _6374_ (.A0(_1471_),
    .A1(_1494_),
    .A2(_1572_),
    .A3(_1580_),
    .S0(net192),
    .S1(net188),
    .X(_3383_));
 sky130_fd_sc_hd__mux2_1 _6375_ (.A0(_3316_),
    .A1(_3383_),
    .S(net198),
    .X(_3384_));
 sky130_fd_sc_hd__mux2_1 _6376_ (.A0(_3251_),
    .A1(_3384_),
    .S(net205),
    .X(_3385_));
 sky130_fd_sc_hd__a2bb2o_1 _6377_ (.A1_N(net180),
    .A2_N(_3385_),
    .B1(_3108_),
    .B2(_2778_),
    .X(_3386_));
 sky130_fd_sc_hd__a21oi_1 _6378_ (.A1(net183),
    .A2(_3113_),
    .B1(_3151_),
    .Y(_3387_));
 sky130_fd_sc_hd__a221o_1 _6379_ (.A1(_1586_),
    .A2(net299),
    .B1(net349),
    .B2(_1584_),
    .C1(net208),
    .X(_3388_));
 sky130_fd_sc_hd__nor2_1 _6380_ (.A(_2765_),
    .B(_3380_),
    .Y(_3389_));
 sky130_fd_sc_hd__a311o_1 _6381_ (.A1(net183),
    .A2(_2931_),
    .A3(_3036_),
    .B1(_3388_),
    .C1(_3389_),
    .X(_3390_));
 sky130_fd_sc_hd__o21ai_1 _6382_ (.A1(net301),
    .A2(_3382_),
    .B1(_3386_),
    .Y(_3391_));
 sky130_fd_sc_hd__a21oi_1 _6383_ (.A1(_1587_),
    .A2(net208),
    .B1(net464),
    .Y(_3392_));
 sky130_fd_sc_hd__o31a_1 _6384_ (.A1(_3387_),
    .A2(_3390_),
    .A3(_3391_),
    .B1(_3392_),
    .X(_0873_));
 sky130_fd_sc_hd__a21oi_2 _6385_ (.A1(_3377_),
    .A2(_3381_),
    .B1(_3378_),
    .Y(_3393_));
 sky130_fd_sc_hd__xnor2_1 _6386_ (.A(_1560_),
    .B(net353),
    .Y(_3394_));
 sky130_fd_sc_hd__and2_1 _6387_ (.A(_1557_),
    .B(_3394_),
    .X(_3395_));
 sky130_fd_sc_hd__or2_1 _6388_ (.A(_1557_),
    .B(_3394_),
    .X(_3396_));
 sky130_fd_sc_hd__and2b_1 _6389_ (.A_N(_3395_),
    .B(_3396_),
    .X(_3397_));
 sky130_fd_sc_hd__xnor2_1 _6390_ (.A(_3393_),
    .B(_3397_),
    .Y(_3398_));
 sky130_fd_sc_hd__nor2_1 _6391_ (.A(net301),
    .B(_3398_),
    .Y(_3399_));
 sky130_fd_sc_hd__mux4_1 _6392_ (.A0(_1494_),
    .A1(_1572_),
    .A2(_1580_),
    .A3(_1557_),
    .S0(net193),
    .S1(net189),
    .X(_3400_));
 sky130_fd_sc_hd__or2_1 _6393_ (.A(net200),
    .B(_3334_),
    .X(_3401_));
 sky130_fd_sc_hd__o21a_1 _6394_ (.A1(net194),
    .A2(_3400_),
    .B1(net204),
    .X(_3402_));
 sky130_fd_sc_hd__a221o_1 _6395_ (.A1(net203),
    .A2(_3265_),
    .B1(_3401_),
    .B2(_3402_),
    .C1(net180),
    .X(_3403_));
 sky130_fd_sc_hd__o211a_1 _6396_ (.A1(net183),
    .A2(_3125_),
    .B1(_3403_),
    .C1(_2775_),
    .X(_3404_));
 sky130_fd_sc_hd__a21oi_1 _6397_ (.A1(_1721_),
    .A2(_3131_),
    .B1(_3151_),
    .Y(_3405_));
 sky130_fd_sc_hd__a221o_1 _6398_ (.A1(_1561_),
    .A2(net300),
    .B1(net349),
    .B2(_1560_),
    .C1(_2772_),
    .X(_3406_));
 sky130_fd_sc_hd__a221o_1 _6399_ (.A1(_1563_),
    .A2(net351),
    .B1(_2958_),
    .B2(_3322_),
    .C1(_3406_),
    .X(_3407_));
 sky130_fd_sc_hd__a21oi_1 _6400_ (.A1(net2387),
    .A2(net208),
    .B1(net464),
    .Y(_3408_));
 sky130_fd_sc_hd__o41a_1 _6401_ (.A1(_3399_),
    .A2(_3404_),
    .A3(_3405_),
    .A4(_3407_),
    .B1(_3408_),
    .X(_0874_));
 sky130_fd_sc_hd__o21ai_1 _6402_ (.A1(_3393_),
    .A2(_3395_),
    .B1(_3396_),
    .Y(_3409_));
 sky130_fd_sc_hd__nor2_1 _6403_ (.A(_1598_),
    .B(_2760_),
    .Y(_3410_));
 sky130_fd_sc_hd__or2_1 _6404_ (.A(_1598_),
    .B(_2760_),
    .X(_3411_));
 sky130_fd_sc_hd__nor2_1 _6405_ (.A(_1599_),
    .B(net353),
    .Y(_3412_));
 sky130_fd_sc_hd__nand2_1 _6406_ (.A(_1598_),
    .B(_2760_),
    .Y(_3413_));
 sky130_fd_sc_hd__o221a_1 _6407_ (.A1(_3393_),
    .A2(_3395_),
    .B1(_3410_),
    .B2(_3412_),
    .C1(_3396_),
    .X(_3414_));
 sky130_fd_sc_hd__a311o_1 _6408_ (.A1(_3409_),
    .A2(_3411_),
    .A3(_3413_),
    .B1(_3414_),
    .C1(net302),
    .X(_3415_));
 sky130_fd_sc_hd__mux4_1 _6409_ (.A0(_1557_),
    .A1(_1572_),
    .A2(_1594_),
    .A3(_1580_),
    .S0(net185),
    .S1(net192),
    .X(_3416_));
 sky130_fd_sc_hd__mux2_1 _6410_ (.A0(_3351_),
    .A1(_3416_),
    .S(net198),
    .X(_3417_));
 sky130_fd_sc_hd__mux2_1 _6411_ (.A0(_3284_),
    .A1(_3417_),
    .S(net205),
    .X(_3418_));
 sky130_fd_sc_hd__mux2_1 _6412_ (.A0(_3146_),
    .A1(_3418_),
    .S(net183),
    .X(_3419_));
 sky130_fd_sc_hd__a221o_1 _6413_ (.A1(_1594_),
    .A2(_2727_),
    .B1(net350),
    .B2(_1592_),
    .C1(net208),
    .X(_3420_));
 sky130_fd_sc_hd__a221o_1 _6414_ (.A1(_1599_),
    .A2(net351),
    .B1(net299),
    .B2(_1597_),
    .C1(_3420_),
    .X(_3421_));
 sky130_fd_sc_hd__a22o_1 _6415_ (.A1(_2983_),
    .A2(_3322_),
    .B1(_3419_),
    .B2(_2775_),
    .X(_3422_));
 sky130_fd_sc_hd__nor2_1 _6416_ (.A(_3421_),
    .B(_3422_),
    .Y(_3423_));
 sky130_fd_sc_hd__a221oi_1 _6417_ (.A1(net2354),
    .A2(net209),
    .B1(_3415_),
    .B2(_3423_),
    .C1(net464),
    .Y(_0875_));
 sky130_fd_sc_hd__and2_1 _6418_ (.A(net455),
    .B(net1342),
    .X(_0876_));
 sky130_fd_sc_hd__and2_1 _6419_ (.A(net455),
    .B(net1716),
    .X(_0877_));
 sky130_fd_sc_hd__and2_1 _6420_ (.A(net455),
    .B(net795),
    .X(_0878_));
 sky130_fd_sc_hd__nor2_2 _6421_ (.A(net468),
    .B(_1678_),
    .Y(_0879_));
 sky130_fd_sc_hd__o31a_2 _6422_ (.A1(_1691_),
    .A2(_1692_),
    .A3(net2307),
    .B1(net458),
    .X(_0880_));
 sky130_fd_sc_hd__nor2_1 _6423_ (.A(net461),
    .B(net2161),
    .Y(_0881_));
 sky130_fd_sc_hd__nor2_1 _6424_ (.A(net466),
    .B(net2193),
    .Y(_0882_));
 sky130_fd_sc_hd__and2_1 _6425_ (.A(net454),
    .B(net2298),
    .X(_0883_));
 sky130_fd_sc_hd__and2_1 _6426_ (.A(net445),
    .B(_1744_),
    .X(_0884_));
 sky130_fd_sc_hd__and2_1 _6427_ (.A(net447),
    .B(net2300),
    .X(_0885_));
 sky130_fd_sc_hd__and2_1 _6428_ (.A(net436),
    .B(net2222),
    .X(_0886_));
 sky130_fd_sc_hd__nor2_1 _6429_ (.A(net466),
    .B(net2296),
    .Y(_0887_));
 sky130_fd_sc_hd__and2_1 _6430_ (.A(net448),
    .B(net2237),
    .X(_0888_));
 sky130_fd_sc_hd__and2_1 _6431_ (.A(net457),
    .B(net2257),
    .X(_0889_));
 sky130_fd_sc_hd__and2_1 _6432_ (.A(net445),
    .B(net2268),
    .X(_0890_));
 sky130_fd_sc_hd__and2_1 _6433_ (.A(net450),
    .B(net2275),
    .X(_0891_));
 sky130_fd_sc_hd__and2_1 _6434_ (.A(net431),
    .B(net2241),
    .X(_0892_));
 sky130_fd_sc_hd__and2_1 _6435_ (.A(net427),
    .B(net2159),
    .X(_0893_));
 sky130_fd_sc_hd__and2_1 _6436_ (.A(net427),
    .B(net2303),
    .X(_0894_));
 sky130_fd_sc_hd__and2_1 _6437_ (.A(net432),
    .B(net2200),
    .X(_0895_));
 sky130_fd_sc_hd__a31oi_1 _6438_ (.A1(_1522_),
    .A2(_1523_),
    .A3(_1524_),
    .B1(net467),
    .Y(_0896_));
 sky130_fd_sc_hd__and2_1 _6439_ (.A(net454),
    .B(net2289),
    .X(_0897_));
 sky130_fd_sc_hd__and2_1 _6440_ (.A(net432),
    .B(net2285),
    .X(_0898_));
 sky130_fd_sc_hd__nor2_2 _6441_ (.A(net461),
    .B(_1616_),
    .Y(_0899_));
 sky130_fd_sc_hd__and2_1 _6442_ (.A(net428),
    .B(net2261),
    .X(_0900_));
 sky130_fd_sc_hd__and2_1 _6443_ (.A(net454),
    .B(net2266),
    .X(_0901_));
 sky130_fd_sc_hd__and2_1 _6444_ (.A(net435),
    .B(_1631_),
    .X(_0902_));
 sky130_fd_sc_hd__nor2_1 _6445_ (.A(net468),
    .B(_1482_),
    .Y(_0903_));
 sky130_fd_sc_hd__and2_1 _6446_ (.A(net439),
    .B(net2293),
    .X(_0904_));
 sky130_fd_sc_hd__and2_1 _6447_ (.A(net435),
    .B(_1473_),
    .X(_0905_));
 sky130_fd_sc_hd__nor2_2 _6448_ (.A(net461),
    .B(_1496_),
    .Y(_0906_));
 sky130_fd_sc_hd__and2_1 _6449_ (.A(net428),
    .B(net2263),
    .X(_0907_));
 sky130_fd_sc_hd__nor2_1 _6450_ (.A(net461),
    .B(net2150),
    .Y(_0908_));
 sky130_fd_sc_hd__and2_1 _6451_ (.A(net441),
    .B(net2281),
    .X(_0909_));
 sky130_fd_sc_hd__and2_1 _6452_ (.A(net435),
    .B(_1591_),
    .X(_0910_));
 sky130_fd_sc_hd__and2_1 _6453_ (.A(net427),
    .B(net1999),
    .X(_0911_));
 sky130_fd_sc_hd__and2_1 _6454_ (.A(net453),
    .B(net2399),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_1 _6455_ (.A0(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .S(net467),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_1 _6456_ (.A0(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .S(net467),
    .X(_0914_));
 sky130_fd_sc_hd__mux2_1 _6457_ (.A0(net2094),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .S(net467),
    .X(_0915_));
 sky130_fd_sc_hd__mux2_1 _6458_ (.A0(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ),
    .A1(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .S(net467),
    .X(_0916_));
 sky130_fd_sc_hd__and2_1 _6459_ (.A(net451),
    .B(net680),
    .X(_0917_));
 sky130_fd_sc_hd__and2_1 _6460_ (.A(net452),
    .B(net799),
    .X(_0918_));
 sky130_fd_sc_hd__and2_1 _6461_ (.A(net441),
    .B(net789),
    .X(_0919_));
 sky130_fd_sc_hd__and2_1 _6462_ (.A(net442),
    .B(net751),
    .X(_0920_));
 sky130_fd_sc_hd__and2_1 _6463_ (.A(net451),
    .B(net797),
    .X(_0921_));
 sky130_fd_sc_hd__and2_1 _6464_ (.A(net452),
    .B(net606),
    .X(_0922_));
 sky130_fd_sc_hd__and2_1 _6465_ (.A(net451),
    .B(net705),
    .X(_0923_));
 sky130_fd_sc_hd__and2_1 _6466_ (.A(net451),
    .B(net688),
    .X(_0924_));
 sky130_fd_sc_hd__and2_1 _6467_ (.A(net455),
    .B(net618),
    .X(_0925_));
 sky130_fd_sc_hd__and2_1 _6468_ (.A(net454),
    .B(net612),
    .X(_0926_));
 sky130_fd_sc_hd__and2_1 _6469_ (.A(net457),
    .B(net674),
    .X(_0927_));
 sky130_fd_sc_hd__and2_1 _6470_ (.A(net456),
    .B(net785),
    .X(_0928_));
 sky130_fd_sc_hd__and2_1 _6471_ (.A(net455),
    .B(net616),
    .X(_0929_));
 sky130_fd_sc_hd__and2_1 _6472_ (.A(net436),
    .B(net644),
    .X(_0930_));
 sky130_fd_sc_hd__and2_1 _6473_ (.A(net435),
    .B(net775),
    .X(_0931_));
 sky130_fd_sc_hd__and2_1 _6474_ (.A(net438),
    .B(net620),
    .X(_0932_));
 sky130_fd_sc_hd__and2_1 _6475_ (.A(net440),
    .B(net739),
    .X(_0933_));
 sky130_fd_sc_hd__and2_1 _6476_ (.A(net437),
    .B(net771),
    .X(_0934_));
 sky130_fd_sc_hd__and2_1 _6477_ (.A(net438),
    .B(net697),
    .X(_0935_));
 sky130_fd_sc_hd__and2_1 _6478_ (.A(net443),
    .B(net841),
    .X(_0936_));
 sky130_fd_sc_hd__and2_1 _6479_ (.A(net438),
    .B(net741),
    .X(_0937_));
 sky130_fd_sc_hd__and2_1 _6480_ (.A(net436),
    .B(net678),
    .X(_0938_));
 sky130_fd_sc_hd__and2_1 _6481_ (.A(net438),
    .B(net636),
    .X(_0939_));
 sky130_fd_sc_hd__and2_1 _6482_ (.A(net440),
    .B(net634),
    .X(_0940_));
 sky130_fd_sc_hd__and2_1 _6483_ (.A(net440),
    .B(net638),
    .X(_0941_));
 sky130_fd_sc_hd__and2_1 _6484_ (.A(net440),
    .B(net763),
    .X(_0942_));
 sky130_fd_sc_hd__and2_1 _6485_ (.A(net441),
    .B(net666),
    .X(_0943_));
 sky130_fd_sc_hd__and2_1 _6486_ (.A(net440),
    .B(net630),
    .X(_0944_));
 sky130_fd_sc_hd__and2_1 _6487_ (.A(net441),
    .B(net765),
    .X(_0945_));
 sky130_fd_sc_hd__and2_1 _6488_ (.A(net441),
    .B(net733),
    .X(_0946_));
 sky130_fd_sc_hd__and2_1 _6489_ (.A(net453),
    .B(net787),
    .X(_0947_));
 sky130_fd_sc_hd__and2_1 _6490_ (.A(net453),
    .B(net761),
    .X(_0948_));
 sky130_fd_sc_hd__and2_1 _6491_ (.A(net451),
    .B(net717),
    .X(_0949_));
 sky130_fd_sc_hd__and2_1 _6492_ (.A(net452),
    .B(net650),
    .X(_0950_));
 sky130_fd_sc_hd__and2_1 _6493_ (.A(net442),
    .B(net745),
    .X(_0951_));
 sky130_fd_sc_hd__and2_1 _6494_ (.A(net452),
    .B(net676),
    .X(_0952_));
 sky130_fd_sc_hd__and2_1 _6495_ (.A(net451),
    .B(net608),
    .X(_0953_));
 sky130_fd_sc_hd__and2_1 _6496_ (.A(net441),
    .B(net737),
    .X(_0954_));
 sky130_fd_sc_hd__and2_1 _6497_ (.A(net451),
    .B(net725),
    .X(_0955_));
 sky130_fd_sc_hd__and2_1 _6498_ (.A(net451),
    .B(net699),
    .X(_0956_));
 sky130_fd_sc_hd__and2_1 _6499_ (.A(net455),
    .B(net773),
    .X(_0957_));
 sky130_fd_sc_hd__and2_1 _6500_ (.A(net453),
    .B(net769),
    .X(_0958_));
 sky130_fd_sc_hd__and2_1 _6501_ (.A(net455),
    .B(net701),
    .X(_0959_));
 sky130_fd_sc_hd__and2_1 _6502_ (.A(net456),
    .B(net614),
    .X(_0960_));
 sky130_fd_sc_hd__and2_1 _6503_ (.A(net456),
    .B(net729),
    .X(_0961_));
 sky130_fd_sc_hd__and2_1 _6504_ (.A(net436),
    .B(net642),
    .X(_0962_));
 sky130_fd_sc_hd__and2_1 _6505_ (.A(net436),
    .B(net662),
    .X(_0963_));
 sky130_fd_sc_hd__and2_1 _6506_ (.A(net438),
    .B(net628),
    .X(_0964_));
 sky130_fd_sc_hd__and2_1 _6507_ (.A(net440),
    .B(net715),
    .X(_0965_));
 sky130_fd_sc_hd__and2_1 _6508_ (.A(net437),
    .B(net624),
    .X(_0966_));
 sky130_fd_sc_hd__and2_1 _6509_ (.A(net438),
    .B(net713),
    .X(_0967_));
 sky130_fd_sc_hd__and2_1 _6510_ (.A(net443),
    .B(net825),
    .X(_0968_));
 sky130_fd_sc_hd__and2_1 _6511_ (.A(net438),
    .B(net626),
    .X(_0969_));
 sky130_fd_sc_hd__and2_1 _6512_ (.A(net436),
    .B(net658),
    .X(_0970_));
 sky130_fd_sc_hd__and2_1 _6513_ (.A(net438),
    .B(net664),
    .X(_0971_));
 sky130_fd_sc_hd__and2_1 _6514_ (.A(net440),
    .B(net652),
    .X(_0972_));
 sky130_fd_sc_hd__and2_1 _6515_ (.A(net439),
    .B(net646),
    .X(_0973_));
 sky130_fd_sc_hd__and2_1 _6516_ (.A(net440),
    .B(net793),
    .X(_0974_));
 sky130_fd_sc_hd__and2_1 _6517_ (.A(net441),
    .B(net692),
    .X(_0975_));
 sky130_fd_sc_hd__and2_1 _6518_ (.A(net440),
    .B(net779),
    .X(_0976_));
 sky130_fd_sc_hd__and2_1 _6519_ (.A(net442),
    .B(net767),
    .X(_0977_));
 sky130_fd_sc_hd__and2_1 _6520_ (.A(net441),
    .B(net686),
    .X(_0978_));
 sky130_fd_sc_hd__and2_1 _6521_ (.A(net457),
    .B(net31),
    .X(_0979_));
 sky130_fd_sc_hd__and2_1 _6522_ (.A(net447),
    .B(net42),
    .X(_0980_));
 sky130_fd_sc_hd__and2_1 _6523_ (.A(net450),
    .B(net53),
    .X(_0981_));
 sky130_fd_sc_hd__and2_1 _6524_ (.A(net440),
    .B(net56),
    .X(_0982_));
 sky130_fd_sc_hd__and2_1 _6525_ (.A(net438),
    .B(net57),
    .X(_0983_));
 sky130_fd_sc_hd__and2_1 _6526_ (.A(net439),
    .B(net58),
    .X(_0984_));
 sky130_fd_sc_hd__and2_1 _6527_ (.A(net444),
    .B(net59),
    .X(_0985_));
 sky130_fd_sc_hd__and2_1 _6528_ (.A(net427),
    .B(net60),
    .X(_0986_));
 sky130_fd_sc_hd__and2_1 _6529_ (.A(net457),
    .B(net61),
    .X(_0987_));
 sky130_fd_sc_hd__and2_1 _6530_ (.A(net429),
    .B(net62),
    .X(_0988_));
 sky130_fd_sc_hd__and2_1 _6531_ (.A(net448),
    .B(net32),
    .X(_0989_));
 sky130_fd_sc_hd__and2_1 _6532_ (.A(net447),
    .B(net33),
    .X(_0990_));
 sky130_fd_sc_hd__and2_1 _6533_ (.A(net456),
    .B(net34),
    .X(_0991_));
 sky130_fd_sc_hd__and2_1 _6534_ (.A(net455),
    .B(net35),
    .X(_0992_));
 sky130_fd_sc_hd__and2_1 _6535_ (.A(net456),
    .B(net36),
    .X(_0993_));
 sky130_fd_sc_hd__and2_1 _6536_ (.A(net435),
    .B(net37),
    .X(_0994_));
 sky130_fd_sc_hd__and2_1 _6537_ (.A(net435),
    .B(net38),
    .X(_0995_));
 sky130_fd_sc_hd__and2_1 _6538_ (.A(net438),
    .B(net39),
    .X(_0996_));
 sky130_fd_sc_hd__and2_1 _6539_ (.A(net442),
    .B(net40),
    .X(_0997_));
 sky130_fd_sc_hd__and2_1 _6540_ (.A(net427),
    .B(net41),
    .X(_0998_));
 sky130_fd_sc_hd__and2_1 _6541_ (.A(net438),
    .B(net43),
    .X(_0999_));
 sky130_fd_sc_hd__and2_1 _6542_ (.A(net450),
    .B(net44),
    .X(_1000_));
 sky130_fd_sc_hd__and2_1 _6543_ (.A(net436),
    .B(net45),
    .X(_1001_));
 sky130_fd_sc_hd__and2_1 _6544_ (.A(net427),
    .B(net46),
    .X(_1002_));
 sky130_fd_sc_hd__and2_1 _6545_ (.A(net436),
    .B(net47),
    .X(_1003_));
 sky130_fd_sc_hd__and2_1 _6546_ (.A(net450),
    .B(net48),
    .X(_1004_));
 sky130_fd_sc_hd__and2_1 _6547_ (.A(net447),
    .B(net49),
    .X(_1005_));
 sky130_fd_sc_hd__and2_1 _6548_ (.A(net456),
    .B(net50),
    .X(_1006_));
 sky130_fd_sc_hd__and2_1 _6549_ (.A(net448),
    .B(net51),
    .X(_1007_));
 sky130_fd_sc_hd__and2_1 _6550_ (.A(net438),
    .B(net52),
    .X(_1008_));
 sky130_fd_sc_hd__and2_1 _6551_ (.A(net439),
    .B(net54),
    .X(_1009_));
 sky130_fd_sc_hd__and2_1 _6552_ (.A(net457),
    .B(net55),
    .X(_1010_));
 sky130_fd_sc_hd__nand2_1 _6553_ (.A(net1988),
    .B(_2687_),
    .Y(_3424_));
 sky130_fd_sc_hd__and4_1 _6554_ (.A(net1989),
    .B(_2711_),
    .C(_2715_),
    .D(_3424_),
    .X(_3425_));
 sky130_fd_sc_hd__a21oi_1 _6555_ (.A1(_2176_),
    .A2(_3425_),
    .B1(net160),
    .Y(_1044_));
 sky130_fd_sc_hd__or3b_4 _6556_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ),
    .C_N(_2653_),
    .X(_3426_));
 sky130_fd_sc_hd__nor2_2 _6557_ (.A(_2655_),
    .B(_3426_),
    .Y(_3427_));
 sky130_fd_sc_hd__or2_1 _6558_ (.A(_2655_),
    .B(_3426_),
    .X(_3428_));
 sky130_fd_sc_hd__nor2_2 _6559_ (.A(net466),
    .B(net297),
    .Y(_3429_));
 sky130_fd_sc_hd__nand2_1 _6560_ (.A(net450),
    .B(_3428_),
    .Y(_3430_));
 sky130_fd_sc_hd__a22o_1 _6561_ (.A1(net356),
    .A2(net298),
    .B1(net252),
    .B2(net1252),
    .X(_1045_));
 sky130_fd_sc_hd__a22o_1 _6562_ (.A1(_1689_),
    .A2(net298),
    .B1(net252),
    .B2(net1328),
    .X(_1046_));
 sky130_fd_sc_hd__o22a_1 _6563_ (.A1(net329),
    .A2(_3428_),
    .B1(_3430_),
    .B2(net909),
    .X(_1047_));
 sky130_fd_sc_hd__o22a_1 _6564_ (.A1(net330),
    .A2(_3428_),
    .B1(_3430_),
    .B2(net885),
    .X(_1048_));
 sky130_fd_sc_hd__a22o_1 _6565_ (.A1(net327),
    .A2(net297),
    .B1(net251),
    .B2(net1668),
    .X(_1049_));
 sky130_fd_sc_hd__a22o_1 _6566_ (.A1(net325),
    .A2(net298),
    .B1(net252),
    .B2(net1700),
    .X(_1050_));
 sky130_fd_sc_hd__a22o_1 _6567_ (.A1(net328),
    .A2(net298),
    .B1(net252),
    .B2(net1546),
    .X(_1051_));
 sky130_fd_sc_hd__a22o_1 _6568_ (.A1(net326),
    .A2(net297),
    .B1(net251),
    .B2(net1334),
    .X(_1052_));
 sky130_fd_sc_hd__a22o_1 _6569_ (.A1(net323),
    .A2(net298),
    .B1(net252),
    .B2(net1009),
    .X(_1053_));
 sky130_fd_sc_hd__a22o_1 _6570_ (.A1(net321),
    .A2(net298),
    .B1(net252),
    .B2(net1670),
    .X(_1054_));
 sky130_fd_sc_hd__a22o_1 _6571_ (.A1(net324),
    .A2(net298),
    .B1(net252),
    .B2(net1442),
    .X(_1055_));
 sky130_fd_sc_hd__a22o_1 _6572_ (.A1(net322),
    .A2(net297),
    .B1(net251),
    .B2(net1456),
    .X(_1056_));
 sky130_fd_sc_hd__a22o_1 _6573_ (.A1(net319),
    .A2(net298),
    .B1(net252),
    .B2(net1542),
    .X(_1057_));
 sky130_fd_sc_hd__a22o_1 _6574_ (.A1(net317),
    .A2(net298),
    .B1(net252),
    .B2(net1750),
    .X(_1058_));
 sky130_fd_sc_hd__a22o_1 _6575_ (.A1(net320),
    .A2(net298),
    .B1(net252),
    .B2(net1286),
    .X(_1059_));
 sky130_fd_sc_hd__a22o_1 _6576_ (.A1(net318),
    .A2(net297),
    .B1(net251),
    .B2(net1620),
    .X(_1060_));
 sky130_fd_sc_hd__a22o_1 _6577_ (.A1(net341),
    .A2(net298),
    .B1(net251),
    .B2(net1448),
    .X(_1061_));
 sky130_fd_sc_hd__a22o_1 _6578_ (.A1(net340),
    .A2(net298),
    .B1(net252),
    .B2(net1586),
    .X(_1062_));
 sky130_fd_sc_hd__a22o_1 _6579_ (.A1(net339),
    .A2(net297),
    .B1(net251),
    .B2(net1592),
    .X(_1063_));
 sky130_fd_sc_hd__a22o_1 _6580_ (.A1(net338),
    .A2(net297),
    .B1(net251),
    .B2(net1656),
    .X(_1064_));
 sky130_fd_sc_hd__a22o_1 _6581_ (.A1(net333),
    .A2(net297),
    .B1(net251),
    .B2(net1632),
    .X(_1065_));
 sky130_fd_sc_hd__a22o_1 _6582_ (.A1(net331),
    .A2(net298),
    .B1(net252),
    .B2(net1548),
    .X(_1066_));
 sky130_fd_sc_hd__a22o_1 _6583_ (.A1(net334),
    .A2(net297),
    .B1(net251),
    .B2(net1708),
    .X(_1067_));
 sky130_fd_sc_hd__a22o_1 _6584_ (.A1(net332),
    .A2(net297),
    .B1(net251),
    .B2(net1474),
    .X(_1068_));
 sky130_fd_sc_hd__a22o_1 _6585_ (.A1(net343),
    .A2(net297),
    .B1(net251),
    .B2(net1596),
    .X(_1069_));
 sky130_fd_sc_hd__a22o_1 _6586_ (.A1(net348),
    .A2(net298),
    .B1(net252),
    .B2(net991),
    .X(_1070_));
 sky130_fd_sc_hd__a22o_1 _6587_ (.A1(net344),
    .A2(net297),
    .B1(net251),
    .B2(net1526),
    .X(_1071_));
 sky130_fd_sc_hd__a22o_1 _6588_ (.A1(net342),
    .A2(net297),
    .B1(net251),
    .B2(net1060),
    .X(_1072_));
 sky130_fd_sc_hd__a22o_1 _6589_ (.A1(net336),
    .A2(net297),
    .B1(net251),
    .B2(net1764),
    .X(_1073_));
 sky130_fd_sc_hd__a22o_1 _6590_ (.A1(net335),
    .A2(net297),
    .B1(net251),
    .B2(net1250),
    .X(_1074_));
 sky130_fd_sc_hd__a22o_1 _6591_ (.A1(net337),
    .A2(net297),
    .B1(net251),
    .B2(net1568),
    .X(_1075_));
 sky130_fd_sc_hd__a22o_1 _6592_ (.A1(_1589_),
    .A2(net298),
    .B1(net252),
    .B2(net1238),
    .X(_1076_));
 sky130_fd_sc_hd__or3b_1 _6593_ (.A(_2693_),
    .B(net1980),
    .C_N(net2127),
    .X(_3431_));
 sky130_fd_sc_hd__a211o_1 _6594_ (.A1(net2048),
    .A2(net2127),
    .B1(_2693_),
    .C1(net1980),
    .X(_3432_));
 sky130_fd_sc_hd__inv_2 _6595_ (.A(_3432_),
    .Y(_3433_));
 sky130_fd_sc_hd__a21oi_1 _6596_ (.A1(_0067_),
    .A2(_2698_),
    .B1(_2708_),
    .Y(_3434_));
 sky130_fd_sc_hd__nor2_1 _6597_ (.A(_1403_),
    .B(_2693_),
    .Y(_3435_));
 sky130_fd_sc_hd__o21a_1 _6598_ (.A1(_3434_),
    .A2(_3435_),
    .B1(_3431_),
    .X(_3436_));
 sky130_fd_sc_hd__o21ai_1 _6599_ (.A1(_3433_),
    .A2(_3436_),
    .B1(_2692_),
    .Y(_3437_));
 sky130_fd_sc_hd__and3_1 _6600_ (.A(_2685_),
    .B(_2706_),
    .C(_3437_),
    .X(_1077_));
 sky130_fd_sc_hd__nor2_1 _6601_ (.A(_2717_),
    .B(_3426_),
    .Y(_3438_));
 sky130_fd_sc_hd__or2_2 _6602_ (.A(_2717_),
    .B(_3426_),
    .X(_3439_));
 sky130_fd_sc_hd__and2_1 _6603_ (.A(net356),
    .B(net296),
    .X(_3440_));
 sky130_fd_sc_hd__a31o_1 _6604_ (.A1(net454),
    .A2(net1722),
    .A3(net294),
    .B1(_3440_),
    .X(_1078_));
 sky130_fd_sc_hd__nor2_1 _6605_ (.A(_1690_),
    .B(net294),
    .Y(_3441_));
 sky130_fd_sc_hd__a31o_1 _6606_ (.A1(net454),
    .A2(net1786),
    .A3(_3439_),
    .B1(_3441_),
    .X(_1079_));
 sky130_fd_sc_hd__or3_1 _6607_ (.A(net467),
    .B(net2100),
    .C(net296),
    .X(_3442_));
 sky130_fd_sc_hd__o21a_1 _6608_ (.A1(net329),
    .A2(net294),
    .B1(_3442_),
    .X(_1080_));
 sky130_fd_sc_hd__and2_1 _6609_ (.A(net330),
    .B(net296),
    .X(_3443_));
 sky130_fd_sc_hd__a31o_1 _6610_ (.A1(net449),
    .A2(net1903),
    .A3(_3439_),
    .B1(_3443_),
    .X(_1081_));
 sky130_fd_sc_hd__and2_1 _6611_ (.A(net327),
    .B(net295),
    .X(_3444_));
 sky130_fd_sc_hd__a31o_1 _6612_ (.A1(net429),
    .A2(net1925),
    .A3(net293),
    .B1(_3444_),
    .X(_1082_));
 sky130_fd_sc_hd__and2_1 _6613_ (.A(net325),
    .B(net296),
    .X(_3445_));
 sky130_fd_sc_hd__a31o_1 _6614_ (.A1(net445),
    .A2(net1927),
    .A3(net294),
    .B1(_3445_),
    .X(_1083_));
 sky130_fd_sc_hd__and2_1 _6615_ (.A(net328),
    .B(net296),
    .X(_3446_));
 sky130_fd_sc_hd__a31o_1 _6616_ (.A1(net447),
    .A2(net1800),
    .A3(net294),
    .B1(_3446_),
    .X(_1084_));
 sky130_fd_sc_hd__and2_1 _6617_ (.A(net326),
    .B(net295),
    .X(_3447_));
 sky130_fd_sc_hd__a31o_1 _6618_ (.A1(net434),
    .A2(net1824),
    .A3(net293),
    .B1(_3447_),
    .X(_1085_));
 sky130_fd_sc_hd__and2_1 _6619_ (.A(net323),
    .B(net296),
    .X(_3448_));
 sky130_fd_sc_hd__a31o_1 _6620_ (.A1(net459),
    .A2(net1684),
    .A3(net294),
    .B1(_3448_),
    .X(_1086_));
 sky130_fd_sc_hd__and2_1 _6621_ (.A(net321),
    .B(net296),
    .X(_3449_));
 sky130_fd_sc_hd__a31o_1 _6622_ (.A1(net448),
    .A2(net1838),
    .A3(net294),
    .B1(_3449_),
    .X(_1087_));
 sky130_fd_sc_hd__and2_1 _6623_ (.A(net324),
    .B(net296),
    .X(_3450_));
 sky130_fd_sc_hd__a31o_1 _6624_ (.A1(net447),
    .A2(net1915),
    .A3(net294),
    .B1(_3450_),
    .X(_1088_));
 sky130_fd_sc_hd__and2_1 _6625_ (.A(net322),
    .B(net295),
    .X(_3451_));
 sky130_fd_sc_hd__a31o_1 _6626_ (.A1(net433),
    .A2(net1862),
    .A3(net293),
    .B1(_3451_),
    .X(_1089_));
 sky130_fd_sc_hd__and2_1 _6627_ (.A(net319),
    .B(net296),
    .X(_3452_));
 sky130_fd_sc_hd__a31o_1 _6628_ (.A1(net449),
    .A2(net1885),
    .A3(net294),
    .B1(_3452_),
    .X(_1090_));
 sky130_fd_sc_hd__and2_1 _6629_ (.A(net317),
    .B(net296),
    .X(_3453_));
 sky130_fd_sc_hd__a31o_1 _6630_ (.A1(net446),
    .A2(net1985),
    .A3(net294),
    .B1(_3453_),
    .X(_1091_));
 sky130_fd_sc_hd__and2_1 _6631_ (.A(net320),
    .B(net296),
    .X(_3454_));
 sky130_fd_sc_hd__a31o_1 _6632_ (.A1(net444),
    .A2(net1780),
    .A3(net294),
    .B1(_3454_),
    .X(_1092_));
 sky130_fd_sc_hd__and2_1 _6633_ (.A(net318),
    .B(net295),
    .X(_3455_));
 sky130_fd_sc_hd__a31o_1 _6634_ (.A1(net433),
    .A2(net1848),
    .A3(net293),
    .B1(_3455_),
    .X(_1093_));
 sky130_fd_sc_hd__and2_1 _6635_ (.A(net341),
    .B(net295),
    .X(_3456_));
 sky130_fd_sc_hd__a31o_1 _6636_ (.A1(net444),
    .A2(net1782),
    .A3(net293),
    .B1(_3456_),
    .X(_1094_));
 sky130_fd_sc_hd__and2_1 _6637_ (.A(net340),
    .B(net296),
    .X(_3457_));
 sky130_fd_sc_hd__a31o_1 _6638_ (.A1(net445),
    .A2(net1909),
    .A3(net294),
    .B1(_3457_),
    .X(_1095_));
 sky130_fd_sc_hd__and2_1 _6639_ (.A(net339),
    .B(net295),
    .X(_3458_));
 sky130_fd_sc_hd__a31o_1 _6640_ (.A1(net428),
    .A2(net1941),
    .A3(net293),
    .B1(_3458_),
    .X(_1096_));
 sky130_fd_sc_hd__and2_1 _6641_ (.A(net338),
    .B(net295),
    .X(_3459_));
 sky130_fd_sc_hd__a31o_1 _6642_ (.A1(net432),
    .A2(net1929),
    .A3(net293),
    .B1(_3459_),
    .X(_1097_));
 sky130_fd_sc_hd__and2_1 _6643_ (.A(net333),
    .B(net295),
    .X(_3460_));
 sky130_fd_sc_hd__a31o_1 _6644_ (.A1(net428),
    .A2(net1856),
    .A3(net293),
    .B1(_3460_),
    .X(_1098_));
 sky130_fd_sc_hd__and2_1 _6645_ (.A(net331),
    .B(net296),
    .X(_3461_));
 sky130_fd_sc_hd__a31o_1 _6646_ (.A1(net444),
    .A2(net1887),
    .A3(net294),
    .B1(_3461_),
    .X(_1099_));
 sky130_fd_sc_hd__and2_1 _6647_ (.A(net334),
    .B(net295),
    .X(_3462_));
 sky130_fd_sc_hd__a31o_1 _6648_ (.A1(net430),
    .A2(net1911),
    .A3(net293),
    .B1(_3462_),
    .X(_1100_));
 sky130_fd_sc_hd__and2_1 _6649_ (.A(net332),
    .B(net295),
    .X(_3463_));
 sky130_fd_sc_hd__a31o_1 _6650_ (.A1(net429),
    .A2(net1939),
    .A3(net293),
    .B1(_3463_),
    .X(_1101_));
 sky130_fd_sc_hd__and2_1 _6651_ (.A(net343),
    .B(net295),
    .X(_3464_));
 sky130_fd_sc_hd__a31o_1 _6652_ (.A1(net435),
    .A2(net1794),
    .A3(net293),
    .B1(_3464_),
    .X(_1102_));
 sky130_fd_sc_hd__and2_1 _6653_ (.A(net348),
    .B(net295),
    .X(_3465_));
 sky130_fd_sc_hd__a31o_1 _6654_ (.A1(net432),
    .A2(net1895),
    .A3(net293),
    .B1(_3465_),
    .X(_1103_));
 sky130_fd_sc_hd__and2_1 _6655_ (.A(net344),
    .B(net295),
    .X(_3466_));
 sky130_fd_sc_hd__a31o_1 _6656_ (.A1(net429),
    .A2(net1901),
    .A3(net293),
    .B1(_3466_),
    .X(_1104_));
 sky130_fd_sc_hd__and2_1 _6657_ (.A(net342),
    .B(net296),
    .X(_3467_));
 sky130_fd_sc_hd__a31o_1 _6658_ (.A1(net429),
    .A2(net1933),
    .A3(net294),
    .B1(_3467_),
    .X(_1105_));
 sky130_fd_sc_hd__and2_1 _6659_ (.A(net336),
    .B(net295),
    .X(_3468_));
 sky130_fd_sc_hd__a31o_1 _6660_ (.A1(net460),
    .A2(net1891),
    .A3(net293),
    .B1(_3468_),
    .X(_1106_));
 sky130_fd_sc_hd__and2_1 _6661_ (.A(net335),
    .B(net296),
    .X(_3469_));
 sky130_fd_sc_hd__a31o_1 _6662_ (.A1(net437),
    .A2(net1868),
    .A3(net294),
    .B1(_3469_),
    .X(_1107_));
 sky130_fd_sc_hd__and2_1 _6663_ (.A(net337),
    .B(net295),
    .X(_3470_));
 sky130_fd_sc_hd__a31o_1 _6664_ (.A1(net434),
    .A2(net1923),
    .A3(net293),
    .B1(_3470_),
    .X(_1108_));
 sky130_fd_sc_hd__and2_1 _6665_ (.A(net357),
    .B(net295),
    .X(_3471_));
 sky130_fd_sc_hd__a31o_1 _6666_ (.A1(net446),
    .A2(net1943),
    .A3(net293),
    .B1(_3471_),
    .X(_1109_));
 sky130_fd_sc_hd__nor2_4 _6667_ (.A(_2670_),
    .B(_2717_),
    .Y(_3472_));
 sky130_fd_sc_hd__or2_1 _6668_ (.A(_2670_),
    .B(_2717_),
    .X(_3473_));
 sky130_fd_sc_hd__nor2_2 _6669_ (.A(net466),
    .B(net292),
    .Y(_3474_));
 sky130_fd_sc_hd__nand2_1 _6670_ (.A(net450),
    .B(_3473_),
    .Y(_3475_));
 sky130_fd_sc_hd__o22a_1 _6671_ (.A1(net356),
    .A2(_3473_),
    .B1(_3475_),
    .B2(net879),
    .X(_1110_));
 sky130_fd_sc_hd__a22o_1 _6672_ (.A1(_1689_),
    .A2(net292),
    .B1(net250),
    .B2(net1074),
    .X(_1111_));
 sky130_fd_sc_hd__o22a_1 _6673_ (.A1(net329),
    .A2(_3473_),
    .B1(_3475_),
    .B2(net857),
    .X(_1112_));
 sky130_fd_sc_hd__a22o_1 _6674_ (.A1(net330),
    .A2(net292),
    .B1(net250),
    .B2(net1134),
    .X(_1113_));
 sky130_fd_sc_hd__a22o_1 _6675_ (.A1(net327),
    .A2(net291),
    .B1(net249),
    .B2(net1296),
    .X(_1114_));
 sky130_fd_sc_hd__a22o_1 _6676_ (.A1(net325),
    .A2(net292),
    .B1(net250),
    .B2(net1362),
    .X(_1115_));
 sky130_fd_sc_hd__a22o_1 _6677_ (.A1(net328),
    .A2(net292),
    .B1(net250),
    .B2(net1022),
    .X(_1116_));
 sky130_fd_sc_hd__a22o_1 _6678_ (.A1(net326),
    .A2(net291),
    .B1(net249),
    .B2(net1530),
    .X(_1117_));
 sky130_fd_sc_hd__a22o_1 _6679_ (.A1(net323),
    .A2(net292),
    .B1(net250),
    .B2(net971),
    .X(_1118_));
 sky130_fd_sc_hd__a22o_1 _6680_ (.A1(net321),
    .A2(net292),
    .B1(net250),
    .B2(net1178),
    .X(_1119_));
 sky130_fd_sc_hd__a22o_1 _6681_ (.A1(net324),
    .A2(net292),
    .B1(net250),
    .B2(net975),
    .X(_1120_));
 sky130_fd_sc_hd__a22o_1 _6682_ (.A1(net322),
    .A2(net291),
    .B1(net249),
    .B2(net1472),
    .X(_1121_));
 sky130_fd_sc_hd__a22o_1 _6683_ (.A1(net319),
    .A2(net292),
    .B1(net250),
    .B2(net947),
    .X(_1122_));
 sky130_fd_sc_hd__a22o_1 _6684_ (.A1(net317),
    .A2(net292),
    .B1(net250),
    .B2(net1056),
    .X(_1123_));
 sky130_fd_sc_hd__a22o_1 _6685_ (.A1(net320),
    .A2(net292),
    .B1(net250),
    .B2(net1064),
    .X(_1124_));
 sky130_fd_sc_hd__a22o_1 _6686_ (.A1(net318),
    .A2(net291),
    .B1(net249),
    .B2(net1510),
    .X(_1125_));
 sky130_fd_sc_hd__a22o_1 _6687_ (.A1(net341),
    .A2(net292),
    .B1(net250),
    .B2(net1312),
    .X(_1126_));
 sky130_fd_sc_hd__a22o_1 _6688_ (.A1(net340),
    .A2(net292),
    .B1(net250),
    .B2(net1460),
    .X(_1127_));
 sky130_fd_sc_hd__a22o_1 _6689_ (.A1(net339),
    .A2(net291),
    .B1(net249),
    .B2(net1444),
    .X(_1128_));
 sky130_fd_sc_hd__a22o_1 _6690_ (.A1(net338),
    .A2(net291),
    .B1(net249),
    .B2(net1192),
    .X(_1129_));
 sky130_fd_sc_hd__a22o_1 _6691_ (.A1(net333),
    .A2(net291),
    .B1(net249),
    .B2(net1080),
    .X(_1130_));
 sky130_fd_sc_hd__a22o_1 _6692_ (.A1(net331),
    .A2(net292),
    .B1(net250),
    .B2(net1290),
    .X(_1131_));
 sky130_fd_sc_hd__a22o_1 _6693_ (.A1(net334),
    .A2(net291),
    .B1(net249),
    .B2(net1236),
    .X(_1132_));
 sky130_fd_sc_hd__a22o_1 _6694_ (.A1(net332),
    .A2(net291),
    .B1(net249),
    .B2(net1132),
    .X(_1133_));
 sky130_fd_sc_hd__a22o_1 _6695_ (.A1(net343),
    .A2(net291),
    .B1(net249),
    .B2(net1066),
    .X(_1134_));
 sky130_fd_sc_hd__a22o_1 _6696_ (.A1(net348),
    .A2(net291),
    .B1(net249),
    .B2(net1408),
    .X(_1135_));
 sky130_fd_sc_hd__a22o_1 _6697_ (.A1(net344),
    .A2(net291),
    .B1(net249),
    .B2(net1176),
    .X(_1136_));
 sky130_fd_sc_hd__a22o_1 _6698_ (.A1(net342),
    .A2(net291),
    .B1(net249),
    .B2(net1576),
    .X(_1137_));
 sky130_fd_sc_hd__a22o_1 _6699_ (.A1(net336),
    .A2(net291),
    .B1(net249),
    .B2(net1174),
    .X(_1138_));
 sky130_fd_sc_hd__a22o_1 _6700_ (.A1(net335),
    .A2(net291),
    .B1(net249),
    .B2(net1624),
    .X(_1139_));
 sky130_fd_sc_hd__a22o_1 _6701_ (.A1(net337),
    .A2(net291),
    .B1(net249),
    .B2(net1658),
    .X(_1140_));
 sky130_fd_sc_hd__a22o_1 _6702_ (.A1(net357),
    .A2(net292),
    .B1(net250),
    .B2(net1446),
    .X(_1141_));
 sky130_fd_sc_hd__nor2_4 _6703_ (.A(_2654_),
    .B(_2717_),
    .Y(_3476_));
 sky130_fd_sc_hd__or2_1 _6704_ (.A(_2654_),
    .B(_2717_),
    .X(_3477_));
 sky130_fd_sc_hd__nor2_2 _6705_ (.A(net466),
    .B(net290),
    .Y(_3478_));
 sky130_fd_sc_hd__nand2_1 _6706_ (.A(net450),
    .B(_3477_),
    .Y(_3479_));
 sky130_fd_sc_hd__a22o_1 _6707_ (.A1(net356),
    .A2(net290),
    .B1(net248),
    .B2(net1372),
    .X(_1142_));
 sky130_fd_sc_hd__o22a_1 _6708_ (.A1(_1689_),
    .A2(_3477_),
    .B1(_3479_),
    .B2(net867),
    .X(_1143_));
 sky130_fd_sc_hd__o22a_1 _6709_ (.A1(net329),
    .A2(_3477_),
    .B1(_3479_),
    .B2(net831),
    .X(_1144_));
 sky130_fd_sc_hd__a22o_1 _6710_ (.A1(net330),
    .A2(net290),
    .B1(net248),
    .B2(net1320),
    .X(_1145_));
 sky130_fd_sc_hd__a22o_1 _6711_ (.A1(net327),
    .A2(net289),
    .B1(net247),
    .B2(net1626),
    .X(_1146_));
 sky130_fd_sc_hd__a22o_1 _6712_ (.A1(net325),
    .A2(net290),
    .B1(net248),
    .B2(net1040),
    .X(_1147_));
 sky130_fd_sc_hd__a22o_1 _6713_ (.A1(net328),
    .A2(net290),
    .B1(net248),
    .B2(net1378),
    .X(_1148_));
 sky130_fd_sc_hd__a22o_1 _6714_ (.A1(net326),
    .A2(net289),
    .B1(net247),
    .B2(net1196),
    .X(_1149_));
 sky130_fd_sc_hd__a22o_1 _6715_ (.A1(net323),
    .A2(net290),
    .B1(net248),
    .B2(net1186),
    .X(_1150_));
 sky130_fd_sc_hd__a22o_1 _6716_ (.A1(net321),
    .A2(net290),
    .B1(net248),
    .B2(net1156),
    .X(_1151_));
 sky130_fd_sc_hd__a22o_1 _6717_ (.A1(net324),
    .A2(net290),
    .B1(net248),
    .B2(net1032),
    .X(_1152_));
 sky130_fd_sc_hd__a22o_1 _6718_ (.A1(net322),
    .A2(net289),
    .B1(net247),
    .B2(net1468),
    .X(_1153_));
 sky130_fd_sc_hd__a22o_1 _6719_ (.A1(net319),
    .A2(net290),
    .B1(net248),
    .B2(net1044),
    .X(_1154_));
 sky130_fd_sc_hd__a22o_1 _6720_ (.A1(net317),
    .A2(net290),
    .B1(net248),
    .B2(net1606),
    .X(_1155_));
 sky130_fd_sc_hd__a22o_1 _6721_ (.A1(net320),
    .A2(net290),
    .B1(net248),
    .B2(net1206),
    .X(_1156_));
 sky130_fd_sc_hd__a22o_1 _6722_ (.A1(net318),
    .A2(net289),
    .B1(net247),
    .B2(net1308),
    .X(_1157_));
 sky130_fd_sc_hd__a22o_1 _6723_ (.A1(net341),
    .A2(net290),
    .B1(net248),
    .B2(net1188),
    .X(_1158_));
 sky130_fd_sc_hd__a22o_1 _6724_ (.A1(net340),
    .A2(net290),
    .B1(net248),
    .B2(net1702),
    .X(_1159_));
 sky130_fd_sc_hd__a22o_1 _6725_ (.A1(net339),
    .A2(net289),
    .B1(net247),
    .B2(net1230),
    .X(_1160_));
 sky130_fd_sc_hd__a22o_1 _6726_ (.A1(net338),
    .A2(net289),
    .B1(net247),
    .B2(net1696),
    .X(_1161_));
 sky130_fd_sc_hd__a22o_1 _6727_ (.A1(net333),
    .A2(net289),
    .B1(net247),
    .B2(net1574),
    .X(_1162_));
 sky130_fd_sc_hd__a22o_1 _6728_ (.A1(net331),
    .A2(net290),
    .B1(net248),
    .B2(net1706),
    .X(_1163_));
 sky130_fd_sc_hd__a22o_1 _6729_ (.A1(net334),
    .A2(net289),
    .B1(net247),
    .B2(net1398),
    .X(_1164_));
 sky130_fd_sc_hd__a22o_1 _6730_ (.A1(net332),
    .A2(net289),
    .B1(net247),
    .B2(net1142),
    .X(_1165_));
 sky130_fd_sc_hd__a22o_1 _6731_ (.A1(net343),
    .A2(net289),
    .B1(net247),
    .B2(net1402),
    .X(_1166_));
 sky130_fd_sc_hd__a22o_1 _6732_ (.A1(net348),
    .A2(net289),
    .B1(net247),
    .B2(net1616),
    .X(_1167_));
 sky130_fd_sc_hd__a22o_1 _6733_ (.A1(net344),
    .A2(net289),
    .B1(net247),
    .B2(net1160),
    .X(_1168_));
 sky130_fd_sc_hd__a22o_1 _6734_ (.A1(net342),
    .A2(net289),
    .B1(net247),
    .B2(net1578),
    .X(_1169_));
 sky130_fd_sc_hd__a22o_1 _6735_ (.A1(net336),
    .A2(net289),
    .B1(net247),
    .B2(net1376),
    .X(_1170_));
 sky130_fd_sc_hd__a22o_1 _6736_ (.A1(net335),
    .A2(net289),
    .B1(net247),
    .B2(net1258),
    .X(_1171_));
 sky130_fd_sc_hd__a22o_1 _6737_ (.A1(net337),
    .A2(net289),
    .B1(net247),
    .B2(net1360),
    .X(_1172_));
 sky130_fd_sc_hd__a22o_1 _6738_ (.A1(net357),
    .A2(net290),
    .B1(net248),
    .B2(net1240),
    .X(_1173_));
 sky130_fd_sc_hd__nor3_1 _6739_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2660_),
    .Y(_3480_));
 sky130_fd_sc_hd__or3_1 _6740_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2660_),
    .X(_3481_));
 sky130_fd_sc_hd__nor2_1 _6741_ (.A(net466),
    .B(net288),
    .Y(_3482_));
 sky130_fd_sc_hd__nand2_1 _6742_ (.A(net454),
    .B(_3481_),
    .Y(_3483_));
 sky130_fd_sc_hd__o22a_1 _6743_ (.A1(net356),
    .A2(_3481_),
    .B1(_3483_),
    .B2(net903),
    .X(_1174_));
 sky130_fd_sc_hd__o22a_1 _6744_ (.A1(_1689_),
    .A2(_3481_),
    .B1(_3483_),
    .B2(net847),
    .X(_1175_));
 sky130_fd_sc_hd__a22o_1 _6745_ (.A1(net329),
    .A2(net288),
    .B1(net246),
    .B2(net1088),
    .X(_1176_));
 sky130_fd_sc_hd__a22o_1 _6746_ (.A1(net330),
    .A2(net288),
    .B1(net246),
    .B2(net1496),
    .X(_1177_));
 sky130_fd_sc_hd__a22o_1 _6747_ (.A1(net327),
    .A2(net287),
    .B1(net245),
    .B2(net1038),
    .X(_1178_));
 sky130_fd_sc_hd__a22o_1 _6748_ (.A1(net325),
    .A2(net288),
    .B1(net246),
    .B2(net1268),
    .X(_1179_));
 sky130_fd_sc_hd__a22o_1 _6749_ (.A1(net328),
    .A2(net288),
    .B1(net246),
    .B2(net1030),
    .X(_1180_));
 sky130_fd_sc_hd__a22o_1 _6750_ (.A1(net326),
    .A2(net287),
    .B1(net245),
    .B2(net1422),
    .X(_1181_));
 sky130_fd_sc_hd__a22o_1 _6751_ (.A1(net323),
    .A2(net288),
    .B1(net246),
    .B2(net1190),
    .X(_1182_));
 sky130_fd_sc_hd__a22o_1 _6752_ (.A1(net321),
    .A2(net288),
    .B1(net246),
    .B2(net1338),
    .X(_1183_));
 sky130_fd_sc_hd__a22o_1 _6753_ (.A1(net324),
    .A2(net288),
    .B1(net246),
    .B2(net1224),
    .X(_1184_));
 sky130_fd_sc_hd__a22o_1 _6754_ (.A1(net322),
    .A2(net287),
    .B1(net245),
    .B2(net1180),
    .X(_1185_));
 sky130_fd_sc_hd__a22o_1 _6755_ (.A1(net319),
    .A2(net288),
    .B1(net246),
    .B2(net1011),
    .X(_1186_));
 sky130_fd_sc_hd__a22o_1 _6756_ (.A1(net317),
    .A2(net288),
    .B1(net246),
    .B2(net1450),
    .X(_1187_));
 sky130_fd_sc_hd__a22o_1 _6757_ (.A1(net320),
    .A2(net288),
    .B1(net246),
    .B2(net1090),
    .X(_1188_));
 sky130_fd_sc_hd__a22o_1 _6758_ (.A1(net318),
    .A2(net287),
    .B1(net245),
    .B2(net1280),
    .X(_1189_));
 sky130_fd_sc_hd__a22o_1 _6759_ (.A1(net341),
    .A2(net287),
    .B1(net245),
    .B2(net1114),
    .X(_1190_));
 sky130_fd_sc_hd__a22o_1 _6760_ (.A1(net340),
    .A2(net288),
    .B1(net246),
    .B2(net1248),
    .X(_1191_));
 sky130_fd_sc_hd__a22o_1 _6761_ (.A1(net339),
    .A2(net287),
    .B1(net245),
    .B2(net1458),
    .X(_1192_));
 sky130_fd_sc_hd__a22o_1 _6762_ (.A1(net338),
    .A2(net287),
    .B1(net245),
    .B2(net1486),
    .X(_1193_));
 sky130_fd_sc_hd__a22o_1 _6763_ (.A1(net333),
    .A2(net287),
    .B1(net245),
    .B2(net983),
    .X(_1194_));
 sky130_fd_sc_hd__a22o_1 _6764_ (.A1(net331),
    .A2(net288),
    .B1(net246),
    .B2(net1050),
    .X(_1195_));
 sky130_fd_sc_hd__a22o_1 _6765_ (.A1(net334),
    .A2(net287),
    .B1(net245),
    .B2(net1262),
    .X(_1196_));
 sky130_fd_sc_hd__a22o_1 _6766_ (.A1(net332),
    .A2(net287),
    .B1(net245),
    .B2(net1204),
    .X(_1197_));
 sky130_fd_sc_hd__a22o_1 _6767_ (.A1(net343),
    .A2(net287),
    .B1(net245),
    .B2(net1544),
    .X(_1198_));
 sky130_fd_sc_hd__a22o_1 _6768_ (.A1(net348),
    .A2(net287),
    .B1(net245),
    .B2(net1082),
    .X(_1199_));
 sky130_fd_sc_hd__a22o_1 _6769_ (.A1(net344),
    .A2(net287),
    .B1(net245),
    .B2(net1538),
    .X(_1200_));
 sky130_fd_sc_hd__a22o_1 _6770_ (.A1(net342),
    .A2(net287),
    .B1(net246),
    .B2(net1400),
    .X(_1201_));
 sky130_fd_sc_hd__a22o_1 _6771_ (.A1(net336),
    .A2(net287),
    .B1(net245),
    .B2(net1404),
    .X(_1202_));
 sky130_fd_sc_hd__a22o_1 _6772_ (.A1(net335),
    .A2(net288),
    .B1(net245),
    .B2(net1664),
    .X(_1203_));
 sky130_fd_sc_hd__a22o_1 _6773_ (.A1(net337),
    .A2(net287),
    .B1(net245),
    .B2(net1672),
    .X(_1204_));
 sky130_fd_sc_hd__a22o_1 _6774_ (.A1(net357),
    .A2(net288),
    .B1(net246),
    .B2(net1222),
    .X(_1205_));
 sky130_fd_sc_hd__nor2_2 _6775_ (.A(_2661_),
    .B(_3426_),
    .Y(_3484_));
 sky130_fd_sc_hd__or2_4 _6776_ (.A(_2661_),
    .B(_3426_),
    .X(_3485_));
 sky130_fd_sc_hd__and2_1 _6777_ (.A(net356),
    .B(net286),
    .X(_3486_));
 sky130_fd_sc_hd__a31o_1 _6778_ (.A1(net450),
    .A2(net1728),
    .A3(net283),
    .B1(_3486_),
    .X(_1206_));
 sky130_fd_sc_hd__nor2_1 _6779_ (.A(_1690_),
    .B(net283),
    .Y(_3487_));
 sky130_fd_sc_hd__a31o_1 _6780_ (.A1(net449),
    .A2(net1726),
    .A3(net283),
    .B1(_3487_),
    .X(_1207_));
 sky130_fd_sc_hd__and2_1 _6781_ (.A(net329),
    .B(net286),
    .X(_3488_));
 sky130_fd_sc_hd__a31o_1 _6782_ (.A1(net450),
    .A2(net1978),
    .A3(net283),
    .B1(_3488_),
    .X(_1208_));
 sky130_fd_sc_hd__or3_1 _6783_ (.A(net467),
    .B(net2119),
    .C(net286),
    .X(_3489_));
 sky130_fd_sc_hd__o21a_1 _6784_ (.A1(net330),
    .A2(net283),
    .B1(_3489_),
    .X(_1209_));
 sky130_fd_sc_hd__and2_1 _6785_ (.A(net327),
    .B(net285),
    .X(_3490_));
 sky130_fd_sc_hd__a31o_1 _6786_ (.A1(net430),
    .A2(net1907),
    .A3(net284),
    .B1(_3490_),
    .X(_1210_));
 sky130_fd_sc_hd__and2_1 _6787_ (.A(_1740_),
    .B(net286),
    .X(_3491_));
 sky130_fd_sc_hd__a31o_1 _6788_ (.A1(net445),
    .A2(net1963),
    .A3(net283),
    .B1(_3491_),
    .X(_1211_));
 sky130_fd_sc_hd__and2_1 _6789_ (.A(net328),
    .B(net286),
    .X(_3492_));
 sky130_fd_sc_hd__a31o_1 _6790_ (.A1(net447),
    .A2(net1953),
    .A3(net283),
    .B1(_3492_),
    .X(_1212_));
 sky130_fd_sc_hd__and2_1 _6791_ (.A(net326),
    .B(net285),
    .X(_3493_));
 sky130_fd_sc_hd__a31o_1 _6792_ (.A1(net434),
    .A2(net1945),
    .A3(net284),
    .B1(_3493_),
    .X(_1213_));
 sky130_fd_sc_hd__and2_1 _6793_ (.A(net323),
    .B(net286),
    .X(_3494_));
 sky130_fd_sc_hd__a31o_1 _6794_ (.A1(net450),
    .A2(net1808),
    .A3(net283),
    .B1(_3494_),
    .X(_1214_));
 sky130_fd_sc_hd__and2_1 _6795_ (.A(net321),
    .B(net286),
    .X(_3495_));
 sky130_fd_sc_hd__a31o_1 _6796_ (.A1(net448),
    .A2(net1967),
    .A3(net283),
    .B1(_3495_),
    .X(_1215_));
 sky130_fd_sc_hd__and2_1 _6797_ (.A(net324),
    .B(net286),
    .X(_3496_));
 sky130_fd_sc_hd__a31o_1 _6798_ (.A1(net447),
    .A2(net1935),
    .A3(net283),
    .B1(_3496_),
    .X(_1216_));
 sky130_fd_sc_hd__and2_1 _6799_ (.A(net322),
    .B(net285),
    .X(_3497_));
 sky130_fd_sc_hd__a31o_1 _6800_ (.A1(net433),
    .A2(net1955),
    .A3(net284),
    .B1(_3497_),
    .X(_1217_));
 sky130_fd_sc_hd__and2_1 _6801_ (.A(net319),
    .B(net286),
    .X(_3498_));
 sky130_fd_sc_hd__a31o_1 _6802_ (.A1(net449),
    .A2(net1850),
    .A3(net283),
    .B1(_3498_),
    .X(_1218_));
 sky130_fd_sc_hd__and2_1 _6803_ (.A(net317),
    .B(net286),
    .X(_3499_));
 sky130_fd_sc_hd__a31o_1 _6804_ (.A1(net446),
    .A2(net1921),
    .A3(_3485_),
    .B1(_3499_),
    .X(_1219_));
 sky130_fd_sc_hd__and2_1 _6805_ (.A(net320),
    .B(net286),
    .X(_3500_));
 sky130_fd_sc_hd__a31o_1 _6806_ (.A1(net444),
    .A2(net1742),
    .A3(net283),
    .B1(_3500_),
    .X(_1220_));
 sky130_fd_sc_hd__and2_1 _6807_ (.A(net318),
    .B(net285),
    .X(_3501_));
 sky130_fd_sc_hd__a31o_1 _6808_ (.A1(net431),
    .A2(net1959),
    .A3(net284),
    .B1(_3501_),
    .X(_1221_));
 sky130_fd_sc_hd__and2_1 _6809_ (.A(net341),
    .B(net285),
    .X(_3502_));
 sky130_fd_sc_hd__a31o_1 _6810_ (.A1(net432),
    .A2(net1949),
    .A3(net284),
    .B1(_3502_),
    .X(_1222_));
 sky130_fd_sc_hd__and2_1 _6811_ (.A(net340),
    .B(net286),
    .X(_3503_));
 sky130_fd_sc_hd__a31o_1 _6812_ (.A1(net448),
    .A2(net1965),
    .A3(net283),
    .B1(_3503_),
    .X(_1223_));
 sky130_fd_sc_hd__and2_1 _6813_ (.A(net339),
    .B(net285),
    .X(_3504_));
 sky130_fd_sc_hd__a31o_1 _6814_ (.A1(net428),
    .A2(net1947),
    .A3(net284),
    .B1(_3504_),
    .X(_1224_));
 sky130_fd_sc_hd__and2_1 _6815_ (.A(_1543_),
    .B(net285),
    .X(_3505_));
 sky130_fd_sc_hd__a31o_1 _6816_ (.A1(net432),
    .A2(net1899),
    .A3(net284),
    .B1(_3505_),
    .X(_1225_));
 sky130_fd_sc_hd__and2_1 _6817_ (.A(net333),
    .B(net285),
    .X(_3506_));
 sky130_fd_sc_hd__a31o_1 _6818_ (.A1(net431),
    .A2(net1874),
    .A3(net284),
    .B1(_3506_),
    .X(_1226_));
 sky130_fd_sc_hd__and2_1 _6819_ (.A(net331),
    .B(net286),
    .X(_3507_));
 sky130_fd_sc_hd__a31o_1 _6820_ (.A1(net444),
    .A2(net1860),
    .A3(net283),
    .B1(_3507_),
    .X(_1227_));
 sky130_fd_sc_hd__and2_1 _6821_ (.A(net334),
    .B(net285),
    .X(_3508_));
 sky130_fd_sc_hd__a31o_1 _6822_ (.A1(net434),
    .A2(net1766),
    .A3(net284),
    .B1(_3508_),
    .X(_1228_));
 sky130_fd_sc_hd__and2_1 _6823_ (.A(net332),
    .B(net285),
    .X(_3509_));
 sky130_fd_sc_hd__a31o_1 _6824_ (.A1(net428),
    .A2(net1774),
    .A3(net284),
    .B1(_3509_),
    .X(_1229_));
 sky130_fd_sc_hd__and2_1 _6825_ (.A(net343),
    .B(net285),
    .X(_3510_));
 sky130_fd_sc_hd__a31o_1 _6826_ (.A1(net430),
    .A2(net1858),
    .A3(net284),
    .B1(_3510_),
    .X(_1230_));
 sky130_fd_sc_hd__and2_1 _6827_ (.A(net348),
    .B(net286),
    .X(_3511_));
 sky130_fd_sc_hd__a31o_1 _6828_ (.A1(net446),
    .A2(net1746),
    .A3(net283),
    .B1(_3511_),
    .X(_1231_));
 sky130_fd_sc_hd__and2_1 _6829_ (.A(net344),
    .B(net285),
    .X(_3512_));
 sky130_fd_sc_hd__a31o_1 _6830_ (.A1(net430),
    .A2(net1937),
    .A3(net284),
    .B1(_3512_),
    .X(_1232_));
 sky130_fd_sc_hd__and2_1 _6831_ (.A(net342),
    .B(net285),
    .X(_3513_));
 sky130_fd_sc_hd__a31o_1 _6832_ (.A1(net430),
    .A2(net1796),
    .A3(net284),
    .B1(_3513_),
    .X(_1233_));
 sky130_fd_sc_hd__and2_1 _6833_ (.A(net336),
    .B(net285),
    .X(_3514_));
 sky130_fd_sc_hd__a31o_1 _6834_ (.A1(net434),
    .A2(net1931),
    .A3(net284),
    .B1(_3514_),
    .X(_1234_));
 sky130_fd_sc_hd__and2_1 _6835_ (.A(net335),
    .B(net285),
    .X(_3515_));
 sky130_fd_sc_hd__a31o_1 _6836_ (.A1(net430),
    .A2(net1951),
    .A3(net284),
    .B1(_3515_),
    .X(_1235_));
 sky130_fd_sc_hd__and2_1 _6837_ (.A(net337),
    .B(net285),
    .X(_3516_));
 sky130_fd_sc_hd__a31o_1 _6838_ (.A1(net433),
    .A2(net1883),
    .A3(net284),
    .B1(_3516_),
    .X(_1236_));
 sky130_fd_sc_hd__and2_1 _6839_ (.A(net357),
    .B(net286),
    .X(_3517_));
 sky130_fd_sc_hd__a31o_1 _6840_ (.A1(net446),
    .A2(net1812),
    .A3(net283),
    .B1(_3517_),
    .X(_1237_));
 sky130_fd_sc_hd__nor3_1 _6841_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2670_),
    .Y(_3518_));
 sky130_fd_sc_hd__or3_4 _6842_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2670_),
    .X(_3519_));
 sky130_fd_sc_hd__or3_1 _6843_ (.A(net467),
    .B(net2134),
    .C(net282),
    .X(_3520_));
 sky130_fd_sc_hd__o21a_1 _6844_ (.A1(net356),
    .A2(net280),
    .B1(_3520_),
    .X(_1268_));
 sky130_fd_sc_hd__nor2_1 _6845_ (.A(_1690_),
    .B(net280),
    .Y(_3521_));
 sky130_fd_sc_hd__a31o_1 _6846_ (.A1(net454),
    .A2(net1760),
    .A3(net280),
    .B1(_3521_),
    .X(_1269_));
 sky130_fd_sc_hd__and2_1 _6847_ (.A(net329),
    .B(net282),
    .X(_3522_));
 sky130_fd_sc_hd__a31o_1 _6848_ (.A1(net449),
    .A2(net1694),
    .A3(net280),
    .B1(_3522_),
    .X(_1270_));
 sky130_fd_sc_hd__and2_1 _6849_ (.A(net330),
    .B(net282),
    .X(_3523_));
 sky130_fd_sc_hd__a31o_1 _6850_ (.A1(net449),
    .A2(net1917),
    .A3(_3519_),
    .B1(_3523_),
    .X(_1271_));
 sky130_fd_sc_hd__and2_1 _6851_ (.A(net327),
    .B(net281),
    .X(_3524_));
 sky130_fd_sc_hd__a31o_1 _6852_ (.A1(net429),
    .A2(net1881),
    .A3(net279),
    .B1(_3524_),
    .X(_1272_));
 sky130_fd_sc_hd__and2_1 _6853_ (.A(net325),
    .B(net282),
    .X(_3525_));
 sky130_fd_sc_hd__a31o_1 _6854_ (.A1(net444),
    .A2(net1740),
    .A3(net280),
    .B1(_3525_),
    .X(_1273_));
 sky130_fd_sc_hd__and2_1 _6855_ (.A(net328),
    .B(net282),
    .X(_3526_));
 sky130_fd_sc_hd__a31o_1 _6856_ (.A1(net447),
    .A2(net1770),
    .A3(net280),
    .B1(_3526_),
    .X(_1274_));
 sky130_fd_sc_hd__and2_1 _6857_ (.A(net326),
    .B(net281),
    .X(_3527_));
 sky130_fd_sc_hd__a31o_1 _6858_ (.A1(net443),
    .A2(net1752),
    .A3(net279),
    .B1(_3527_),
    .X(_1275_));
 sky130_fd_sc_hd__and2_1 _6859_ (.A(net323),
    .B(net282),
    .X(_3528_));
 sky130_fd_sc_hd__a31o_1 _6860_ (.A1(net453),
    .A2(net1854),
    .A3(net280),
    .B1(_3528_),
    .X(_1276_));
 sky130_fd_sc_hd__and2_1 _6861_ (.A(net321),
    .B(net282),
    .X(_3529_));
 sky130_fd_sc_hd__a31o_1 _6862_ (.A1(net448),
    .A2(net1788),
    .A3(net280),
    .B1(_3529_),
    .X(_1277_));
 sky130_fd_sc_hd__and2_1 _6863_ (.A(net324),
    .B(net282),
    .X(_3530_));
 sky130_fd_sc_hd__a31o_1 _6864_ (.A1(net447),
    .A2(net1826),
    .A3(_3519_),
    .B1(_3530_),
    .X(_1278_));
 sky130_fd_sc_hd__and2_1 _6865_ (.A(net322),
    .B(net281),
    .X(_3531_));
 sky130_fd_sc_hd__a31o_1 _6866_ (.A1(net433),
    .A2(net1768),
    .A3(net279),
    .B1(_3531_),
    .X(_1279_));
 sky130_fd_sc_hd__and2_1 _6867_ (.A(net319),
    .B(net282),
    .X(_3532_));
 sky130_fd_sc_hd__a31o_1 _6868_ (.A1(net449),
    .A2(net1804),
    .A3(net280),
    .B1(_3532_),
    .X(_1280_));
 sky130_fd_sc_hd__and2_1 _6869_ (.A(net317),
    .B(net282),
    .X(_3533_));
 sky130_fd_sc_hd__a31o_1 _6870_ (.A1(net446),
    .A2(net1778),
    .A3(net280),
    .B1(_3533_),
    .X(_1281_));
 sky130_fd_sc_hd__and2_1 _6871_ (.A(net320),
    .B(net282),
    .X(_3534_));
 sky130_fd_sc_hd__a31o_1 _6872_ (.A1(net444),
    .A2(net1720),
    .A3(net280),
    .B1(_3534_),
    .X(_1282_));
 sky130_fd_sc_hd__and2_1 _6873_ (.A(net318),
    .B(net281),
    .X(_3535_));
 sky130_fd_sc_hd__a31o_1 _6874_ (.A1(net428),
    .A2(net1844),
    .A3(net279),
    .B1(_3535_),
    .X(_1283_));
 sky130_fd_sc_hd__and2_1 _6875_ (.A(net341),
    .B(net281),
    .X(_3536_));
 sky130_fd_sc_hd__a31o_1 _6876_ (.A1(net432),
    .A2(net1748),
    .A3(net279),
    .B1(_3536_),
    .X(_1284_));
 sky130_fd_sc_hd__and2_1 _6877_ (.A(net340),
    .B(net282),
    .X(_3537_));
 sky130_fd_sc_hd__a31o_1 _6878_ (.A1(net459),
    .A2(net1976),
    .A3(net280),
    .B1(_3537_),
    .X(_1285_));
 sky130_fd_sc_hd__and2_1 _6879_ (.A(net339),
    .B(net281),
    .X(_3538_));
 sky130_fd_sc_hd__a31o_1 _6880_ (.A1(net428),
    .A2(net1830),
    .A3(net279),
    .B1(_3538_),
    .X(_1286_));
 sky130_fd_sc_hd__and2_1 _6881_ (.A(net338),
    .B(net281),
    .X(_3539_));
 sky130_fd_sc_hd__a31o_1 _6882_ (.A1(net432),
    .A2(net1762),
    .A3(net279),
    .B1(_3539_),
    .X(_1287_));
 sky130_fd_sc_hd__and2_1 _6883_ (.A(net333),
    .B(net281),
    .X(_3540_));
 sky130_fd_sc_hd__a31o_1 _6884_ (.A1(net427),
    .A2(net1798),
    .A3(net279),
    .B1(_3540_),
    .X(_1288_));
 sky130_fd_sc_hd__and2_1 _6885_ (.A(net331),
    .B(net282),
    .X(_3541_));
 sky130_fd_sc_hd__a31o_1 _6886_ (.A1(net444),
    .A2(net1864),
    .A3(net280),
    .B1(_3541_),
    .X(_1289_));
 sky130_fd_sc_hd__and2_1 _6887_ (.A(net334),
    .B(net281),
    .X(_3542_));
 sky130_fd_sc_hd__a31o_1 _6888_ (.A1(net434),
    .A2(net1814),
    .A3(net279),
    .B1(_3542_),
    .X(_1290_));
 sky130_fd_sc_hd__and2_1 _6889_ (.A(net332),
    .B(net281),
    .X(_3543_));
 sky130_fd_sc_hd__a31o_1 _6890_ (.A1(net429),
    .A2(net1732),
    .A3(net279),
    .B1(_3543_),
    .X(_1291_));
 sky130_fd_sc_hd__and2_1 _6891_ (.A(net343),
    .B(net281),
    .X(_3544_));
 sky130_fd_sc_hd__a31o_1 _6892_ (.A1(net435),
    .A2(net1842),
    .A3(net279),
    .B1(_3544_),
    .X(_1292_));
 sky130_fd_sc_hd__and2_1 _6893_ (.A(net348),
    .B(net281),
    .X(_3545_));
 sky130_fd_sc_hd__a31o_1 _6894_ (.A1(net444),
    .A2(net1738),
    .A3(net279),
    .B1(_3545_),
    .X(_1293_));
 sky130_fd_sc_hd__and2_1 _6895_ (.A(net344),
    .B(net281),
    .X(_3546_));
 sky130_fd_sc_hd__a31o_1 _6896_ (.A1(net429),
    .A2(net1870),
    .A3(net280),
    .B1(_3546_),
    .X(_1294_));
 sky130_fd_sc_hd__and2_1 _6897_ (.A(net342),
    .B(net282),
    .X(_3547_));
 sky130_fd_sc_hd__a31o_1 _6898_ (.A1(net430),
    .A2(net1802),
    .A3(net279),
    .B1(_3547_),
    .X(_1295_));
 sky130_fd_sc_hd__and2_1 _6899_ (.A(net336),
    .B(net281),
    .X(_3548_));
 sky130_fd_sc_hd__a31o_1 _6900_ (.A1(net433),
    .A2(net1822),
    .A3(net279),
    .B1(_3548_),
    .X(_1296_));
 sky130_fd_sc_hd__and2_1 _6901_ (.A(net335),
    .B(net282),
    .X(_3549_));
 sky130_fd_sc_hd__a31o_1 _6902_ (.A1(net437),
    .A2(net1714),
    .A3(net280),
    .B1(_3549_),
    .X(_1297_));
 sky130_fd_sc_hd__and2_1 _6903_ (.A(net337),
    .B(net281),
    .X(_3550_));
 sky130_fd_sc_hd__a31o_1 _6904_ (.A1(net431),
    .A2(net1836),
    .A3(net279),
    .B1(_3550_),
    .X(_1298_));
 sky130_fd_sc_hd__and2_1 _6905_ (.A(net357),
    .B(net281),
    .X(_3551_));
 sky130_fd_sc_hd__a31o_1 _6906_ (.A1(net434),
    .A2(net1840),
    .A3(net279),
    .B1(_3551_),
    .X(_1299_));
 sky130_fd_sc_hd__nor3_4 _6907_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2654_),
    .Y(_3552_));
 sky130_fd_sc_hd__or3_4 _6908_ (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ),
    .B(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ),
    .C(_2654_),
    .X(_3553_));
 sky130_fd_sc_hd__and2_1 _6909_ (.A(_1676_),
    .B(net278),
    .X(_3554_));
 sky130_fd_sc_hd__a31o_1 _6910_ (.A1(net454),
    .A2(net1704),
    .A3(net276),
    .B1(_3554_),
    .X(_1300_));
 sky130_fd_sc_hd__or3_1 _6911_ (.A(net467),
    .B(net2123),
    .C(net278),
    .X(_3555_));
 sky130_fd_sc_hd__o21a_1 _6912_ (.A1(_1689_),
    .A2(net276),
    .B1(_3555_),
    .X(_1301_));
 sky130_fd_sc_hd__and2_1 _6913_ (.A(_1665_),
    .B(net278),
    .X(_3556_));
 sky130_fd_sc_hd__a31o_1 _6914_ (.A1(net449),
    .A2(net1734),
    .A3(net276),
    .B1(_3556_),
    .X(_1302_));
 sky130_fd_sc_hd__and2_1 _6915_ (.A(_1652_),
    .B(net278),
    .X(_3557_));
 sky130_fd_sc_hd__a31o_1 _6916_ (.A1(net449),
    .A2(net1818),
    .A3(net276),
    .B1(_3557_),
    .X(_1303_));
 sky130_fd_sc_hd__and2_1 _6917_ (.A(net327),
    .B(net277),
    .X(_3558_));
 sky130_fd_sc_hd__a31o_1 _6918_ (.A1(net429),
    .A2(net1810),
    .A3(net275),
    .B1(_3558_),
    .X(_1304_));
 sky130_fd_sc_hd__and2_1 _6919_ (.A(net2168),
    .B(net276),
    .X(_3559_));
 sky130_fd_sc_hd__a22o_1 _6920_ (.A1(net325),
    .A2(net278),
    .B1(_3559_),
    .B2(net445),
    .X(_1305_));
 sky130_fd_sc_hd__and2_1 _6921_ (.A(net328),
    .B(net278),
    .X(_3560_));
 sky130_fd_sc_hd__a31o_1 _6922_ (.A1(net447),
    .A2(net1744),
    .A3(net276),
    .B1(_3560_),
    .X(_1306_));
 sky130_fd_sc_hd__and2_1 _6923_ (.A(net326),
    .B(net277),
    .X(_3561_));
 sky130_fd_sc_hd__a31o_1 _6924_ (.A1(net434),
    .A2(net1718),
    .A3(net275),
    .B1(_3561_),
    .X(_1307_));
 sky130_fd_sc_hd__and2_1 _6925_ (.A(net323),
    .B(net278),
    .X(_3562_));
 sky130_fd_sc_hd__a31o_1 _6926_ (.A1(net453),
    .A2(net1736),
    .A3(net276),
    .B1(_3562_),
    .X(_1308_));
 sky130_fd_sc_hd__and2_1 _6927_ (.A(net321),
    .B(net278),
    .X(_3563_));
 sky130_fd_sc_hd__a31o_1 _6928_ (.A1(net448),
    .A2(net1756),
    .A3(net276),
    .B1(_3563_),
    .X(_1309_));
 sky130_fd_sc_hd__and2_1 _6929_ (.A(net324),
    .B(net278),
    .X(_3564_));
 sky130_fd_sc_hd__a31o_1 _6930_ (.A1(net447),
    .A2(net1876),
    .A3(net276),
    .B1(_3564_),
    .X(_1310_));
 sky130_fd_sc_hd__and2_1 _6931_ (.A(net322),
    .B(net277),
    .X(_3565_));
 sky130_fd_sc_hd__a31o_1 _6932_ (.A1(net433),
    .A2(net1790),
    .A3(net275),
    .B1(_3565_),
    .X(_1311_));
 sky130_fd_sc_hd__and2_1 _6933_ (.A(net319),
    .B(net278),
    .X(_3566_));
 sky130_fd_sc_hd__a31o_1 _6934_ (.A1(net448),
    .A2(net1828),
    .A3(net276),
    .B1(_3566_),
    .X(_1312_));
 sky130_fd_sc_hd__and2_1 _6935_ (.A(net317),
    .B(net278),
    .X(_3567_));
 sky130_fd_sc_hd__a31o_1 _6936_ (.A1(net446),
    .A2(net1872),
    .A3(net276),
    .B1(_3567_),
    .X(_1313_));
 sky130_fd_sc_hd__and2_1 _6937_ (.A(net320),
    .B(net278),
    .X(_3568_));
 sky130_fd_sc_hd__a31o_1 _6938_ (.A1(net444),
    .A2(net1905),
    .A3(net276),
    .B1(_3568_),
    .X(_1314_));
 sky130_fd_sc_hd__and2_1 _6939_ (.A(net318),
    .B(net277),
    .X(_3569_));
 sky130_fd_sc_hd__a31o_1 _6940_ (.A1(net431),
    .A2(net1834),
    .A3(net275),
    .B1(_3569_),
    .X(_1315_));
 sky130_fd_sc_hd__and2_1 _6941_ (.A(net341),
    .B(net277),
    .X(_3570_));
 sky130_fd_sc_hd__a31o_1 _6942_ (.A1(net432),
    .A2(net1852),
    .A3(net275),
    .B1(_3570_),
    .X(_1316_));
 sky130_fd_sc_hd__and2_1 _6943_ (.A(net2155),
    .B(net276),
    .X(_3571_));
 sky130_fd_sc_hd__a22o_1 _6944_ (.A1(net340),
    .A2(net278),
    .B1(net2156),
    .B2(net445),
    .X(_1317_));
 sky130_fd_sc_hd__and2_1 _6945_ (.A(net339),
    .B(net277),
    .X(_3572_));
 sky130_fd_sc_hd__a31o_1 _6946_ (.A1(net428),
    .A2(net1846),
    .A3(net275),
    .B1(_3572_),
    .X(_1318_));
 sky130_fd_sc_hd__and2_1 _6947_ (.A(net338),
    .B(net277),
    .X(_3573_));
 sky130_fd_sc_hd__a31o_1 _6948_ (.A1(net432),
    .A2(net1974),
    .A3(net275),
    .B1(_3573_),
    .X(_1319_));
 sky130_fd_sc_hd__and2_1 _6949_ (.A(net333),
    .B(net277),
    .X(_3574_));
 sky130_fd_sc_hd__a31o_1 _6950_ (.A1(net427),
    .A2(net1730),
    .A3(net275),
    .B1(_3574_),
    .X(_1320_));
 sky130_fd_sc_hd__and2_1 _6951_ (.A(net331),
    .B(net278),
    .X(_3575_));
 sky130_fd_sc_hd__a31o_1 _6952_ (.A1(net444),
    .A2(net1724),
    .A3(net276),
    .B1(_3575_),
    .X(_1321_));
 sky130_fd_sc_hd__and2_1 _6953_ (.A(net334),
    .B(net277),
    .X(_3576_));
 sky130_fd_sc_hd__a31o_1 _6954_ (.A1(net434),
    .A2(net1832),
    .A3(net275),
    .B1(_3576_),
    .X(_1322_));
 sky130_fd_sc_hd__and2_1 _6955_ (.A(net332),
    .B(net277),
    .X(_3577_));
 sky130_fd_sc_hd__a31o_1 _6956_ (.A1(net427),
    .A2(net1913),
    .A3(net275),
    .B1(_3577_),
    .X(_1323_));
 sky130_fd_sc_hd__and2_1 _6957_ (.A(_1480_),
    .B(net277),
    .X(_3578_));
 sky130_fd_sc_hd__a31o_1 _6958_ (.A1(net435),
    .A2(net1806),
    .A3(net275),
    .B1(_3578_),
    .X(_1324_));
 sky130_fd_sc_hd__and2_1 _6959_ (.A(net348),
    .B(net277),
    .X(_3579_));
 sky130_fd_sc_hd__a31o_1 _6960_ (.A1(net433),
    .A2(net1889),
    .A3(net275),
    .B1(_3579_),
    .X(_1325_));
 sky130_fd_sc_hd__and2_1 _6961_ (.A(net344),
    .B(net277),
    .X(_3580_));
 sky130_fd_sc_hd__a31o_1 _6962_ (.A1(net429),
    .A2(net1754),
    .A3(net275),
    .B1(_3580_),
    .X(_1326_));
 sky130_fd_sc_hd__and2_1 _6963_ (.A(net342),
    .B(net278),
    .X(_3581_));
 sky130_fd_sc_hd__a31o_1 _6964_ (.A1(net429),
    .A2(net1919),
    .A3(net276),
    .B1(_3581_),
    .X(_1327_));
 sky130_fd_sc_hd__and2_1 _6965_ (.A(net336),
    .B(net277),
    .X(_3582_));
 sky130_fd_sc_hd__a31o_1 _6966_ (.A1(net432),
    .A2(net1961),
    .A3(net275),
    .B1(_3582_),
    .X(_1328_));
 sky130_fd_sc_hd__and2_1 _6967_ (.A(net335),
    .B(net277),
    .X(_3583_));
 sky130_fd_sc_hd__a31o_1 _6968_ (.A1(net437),
    .A2(net1776),
    .A3(net275),
    .B1(_3583_),
    .X(_1329_));
 sky130_fd_sc_hd__and2_1 _6969_ (.A(net337),
    .B(net277),
    .X(_3584_));
 sky130_fd_sc_hd__a31o_1 _6970_ (.A1(net431),
    .A2(net1866),
    .A3(net275),
    .B1(_3584_),
    .X(_1330_));
 sky130_fd_sc_hd__and2_1 _6971_ (.A(net357),
    .B(_3552_),
    .X(_3585_));
 sky130_fd_sc_hd__a31o_1 _6972_ (.A1(net446),
    .A2(net1816),
    .A3(_3553_),
    .B1(_3585_),
    .X(_1331_));
 sky130_fd_sc_hd__nor3_1 _6973_ (.A(net160),
    .B(_2688_),
    .C(_2716_),
    .Y(_1332_));
 sky130_fd_sc_hd__or2_1 _6974_ (.A(_2681_),
    .B(_2705_),
    .X(_3586_));
 sky130_fd_sc_hd__and3_1 _6975_ (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .B(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .C(_2701_),
    .X(_3587_));
 sky130_fd_sc_hd__nor2_1 _6976_ (.A(_2697_),
    .B(_3587_),
    .Y(_3588_));
 sky130_fd_sc_hd__and4b_1 _6977_ (.A_N(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .B(_1403_),
    .C(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ),
    .D(_2703_),
    .X(_3589_));
 sky130_fd_sc_hd__a221o_1 _6978_ (.A1(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .A2(_3587_),
    .B1(_3588_),
    .B2(_0064_),
    .C1(_3589_),
    .X(_3590_));
 sky130_fd_sc_hd__o22a_1 _6979_ (.A1(_1403_),
    .A2(_2693_),
    .B1(_2704_),
    .B2(_2681_),
    .X(_3591_));
 sky130_fd_sc_hd__a2bb2o_1 _6980_ (.A1_N(_2693_),
    .A2_N(_2695_),
    .B1(_3590_),
    .B2(_3591_),
    .X(_3592_));
 sky130_fd_sc_hd__nand2_1 _6981_ (.A(_2684_),
    .B(_2705_),
    .Y(_3593_));
 sky130_fd_sc_hd__a31o_1 _6982_ (.A1(_2692_),
    .A2(_3432_),
    .A3(_3592_),
    .B1(_3593_),
    .X(_3594_));
 sky130_fd_sc_hd__and2b_1 _6983_ (.A_N(_3594_),
    .B(_2696_),
    .X(_3595_));
 sky130_fd_sc_hd__mux2_1 _6984_ (.A0(net2048),
    .A1(_3595_),
    .S(_3586_),
    .X(_3596_));
 sky130_fd_sc_hd__nor2_1 _6985_ (.A(net160),
    .B(_3596_),
    .Y(_1333_));
 sky130_fd_sc_hd__nand2b_1 _6986_ (.A_N(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ),
    .B(net2291),
    .Y(_3597_));
 sky130_fd_sc_hd__a22o_1 _6987_ (.A1(_0065_),
    .A2(_3588_),
    .B1(_3597_),
    .B2(_2708_),
    .X(_3598_));
 sky130_fd_sc_hd__a221o_1 _6988_ (.A1(net1980),
    .A2(_2690_),
    .B1(_2693_),
    .B2(_3598_),
    .C1(_3433_),
    .X(_3599_));
 sky130_fd_sc_hd__a21oi_1 _6989_ (.A1(_2691_),
    .A2(_3599_),
    .B1(_3593_),
    .Y(_3600_));
 sky130_fd_sc_hd__mux2_1 _6990_ (.A0(net2048),
    .A1(_3600_),
    .S(_3586_),
    .X(_3601_));
 sky130_fd_sc_hd__nor2_1 _6991_ (.A(net160),
    .B(_3601_),
    .Y(_1334_));
 sky130_fd_sc_hd__a21o_1 _6992_ (.A1(_0066_),
    .A2(_2698_),
    .B1(_3587_),
    .X(_3602_));
 sky130_fd_sc_hd__o31a_1 _6993_ (.A1(net2145),
    .A2(net1980),
    .A3(_2704_),
    .B1(_3602_),
    .X(_3603_));
 sky130_fd_sc_hd__a2bb2o_1 _6994_ (.A1_N(net2048),
    .A2_N(_3431_),
    .B1(_3603_),
    .B2(_2707_),
    .X(_3604_));
 sky130_fd_sc_hd__a21boi_1 _6995_ (.A1(_2694_),
    .A2(_3604_),
    .B1_N(_2696_),
    .Y(_3605_));
 sky130_fd_sc_hd__o21ai_1 _6996_ (.A1(_3593_),
    .A2(_3605_),
    .B1(_3586_),
    .Y(_3606_));
 sky130_fd_sc_hd__o211a_1 _6997_ (.A1(net2048),
    .A2(_3586_),
    .B1(_3606_),
    .C1(_2679_),
    .X(_1335_));
 sky130_fd_sc_hd__and2_1 _6998_ (.A(net454),
    .B(net1614),
    .X(_1336_));
 sky130_fd_sc_hd__and2_1 _6999_ (.A(net454),
    .B(net1498),
    .X(_1337_));
 sky130_fd_sc_hd__and2_1 _7000_ (.A(net449),
    .B(net1184),
    .X(_1338_));
 sky130_fd_sc_hd__and2_1 _7001_ (.A(net449),
    .B(net1686),
    .X(_1339_));
 sky130_fd_sc_hd__and2_1 _7002_ (.A(net429),
    .B(net1326),
    .X(_1340_));
 sky130_fd_sc_hd__and2_1 _7003_ (.A(net444),
    .B(net1652),
    .X(_1341_));
 sky130_fd_sc_hd__and2_1 _7004_ (.A(net447),
    .B(net1302),
    .X(_1342_));
 sky130_fd_sc_hd__and2_1 _7005_ (.A(net443),
    .B(net1292),
    .X(_1343_));
 sky130_fd_sc_hd__and2_1 _7006_ (.A(net453),
    .B(net1336),
    .X(_1344_));
 sky130_fd_sc_hd__and2_1 _7007_ (.A(net448),
    .B(net1676),
    .X(_1345_));
 sky130_fd_sc_hd__and2_1 _7008_ (.A(net447),
    .B(net1324),
    .X(_1346_));
 sky130_fd_sc_hd__and2_1 _7009_ (.A(net433),
    .B(net1610),
    .X(_1347_));
 sky130_fd_sc_hd__and2_1 _7010_ (.A(net449),
    .B(net1556),
    .X(_1348_));
 sky130_fd_sc_hd__and2_1 _7011_ (.A(net446),
    .B(net1482),
    .X(_1349_));
 sky130_fd_sc_hd__and2_1 _7012_ (.A(net444),
    .B(net1348),
    .X(_1350_));
 sky130_fd_sc_hd__and2_1 _7013_ (.A(net428),
    .B(net1598),
    .X(_1351_));
 sky130_fd_sc_hd__and2_1 _7014_ (.A(net432),
    .B(net1432),
    .X(_1352_));
 sky130_fd_sc_hd__and2_1 _7015_ (.A(net445),
    .B(net1648),
    .X(_1353_));
 sky130_fd_sc_hd__and2_1 _7016_ (.A(net428),
    .B(net1518),
    .X(_1354_));
 sky130_fd_sc_hd__and2_1 _7017_ (.A(net432),
    .B(net1612),
    .X(_1355_));
 sky130_fd_sc_hd__and2_1 _7018_ (.A(net427),
    .B(net1636),
    .X(_1356_));
 sky130_fd_sc_hd__and2_1 _7019_ (.A(net444),
    .B(net1628),
    .X(_1357_));
 sky130_fd_sc_hd__and2_1 _7020_ (.A(net434),
    .B(net1514),
    .X(_1358_));
 sky130_fd_sc_hd__and2_1 _7021_ (.A(net429),
    .B(net1346),
    .X(_1359_));
 sky130_fd_sc_hd__and2_1 _7022_ (.A(net435),
    .B(net1692),
    .X(_1360_));
 sky130_fd_sc_hd__and2_1 _7023_ (.A(net433),
    .B(net1540),
    .X(_1361_));
 sky130_fd_sc_hd__and2_1 _7024_ (.A(net429),
    .B(net1452),
    .X(_1362_));
 sky130_fd_sc_hd__and2_1 _7025_ (.A(net430),
    .B(net1618),
    .X(_1363_));
 sky130_fd_sc_hd__and2_1 _7026_ (.A(net434),
    .B(net1674),
    .X(_1364_));
 sky130_fd_sc_hd__and2_1 _7027_ (.A(net437),
    .B(net1500),
    .X(_1365_));
 sky130_fd_sc_hd__and2_1 _7028_ (.A(net428),
    .B(net1508),
    .X(_1366_));
 sky130_fd_sc_hd__and2_1 _7029_ (.A(net446),
    .B(net1588),
    .X(_1367_));
 sky130_fd_sc_hd__and3_1 _7030_ (.A(net2090),
    .B(net173),
    .C(net221),
    .X(_1368_));
 sky130_fd_sc_hd__nand2_4 _7031_ (.A(net2090),
    .B(net1989),
    .Y(_3607_));
 sky130_fd_sc_hd__nand2_1 _7032_ (.A(net2048),
    .B(_2700_),
    .Y(_3608_));
 sky130_fd_sc_hd__a21oi_1 _7033_ (.A1(_3607_),
    .A2(net2049),
    .B1(net159),
    .Y(_1369_));
 sky130_fd_sc_hd__nand2_1 _7034_ (.A(net1971),
    .B(_2700_),
    .Y(_3609_));
 sky130_fd_sc_hd__a21oi_1 _7035_ (.A1(_3607_),
    .A2(net1972),
    .B1(net159),
    .Y(_1370_));
 sky130_fd_sc_hd__nand2_1 _7036_ (.A(net2175),
    .B(_2700_),
    .Y(_3610_));
 sky130_fd_sc_hd__a21oi_1 _7037_ (.A1(_3607_),
    .A2(net2176),
    .B1(net159),
    .Y(_1371_));
 sky130_fd_sc_hd__nand2_1 _7038_ (.A(net1878),
    .B(_2700_),
    .Y(_3611_));
 sky130_fd_sc_hd__a21oi_1 _7039_ (.A1(_3607_),
    .A2(net1879),
    .B1(net159),
    .Y(_1372_));
 sky130_fd_sc_hd__nand2_1 _7040_ (.A(net2188),
    .B(_2700_),
    .Y(_3612_));
 sky130_fd_sc_hd__a21oi_1 _7041_ (.A1(_3607_),
    .A2(net2189),
    .B1(net159),
    .Y(_1373_));
 sky130_fd_sc_hd__nand2_1 _7042_ (.A(net2083),
    .B(_2700_),
    .Y(_3613_));
 sky130_fd_sc_hd__a21oi_1 _7043_ (.A1(_3607_),
    .A2(net2084),
    .B1(net159),
    .Y(_1374_));
 sky130_fd_sc_hd__nand2_1 _7044_ (.A(net2109),
    .B(_2700_),
    .Y(_3614_));
 sky130_fd_sc_hd__a21oi_1 _7045_ (.A1(_3607_),
    .A2(net2110),
    .B1(net159),
    .Y(_1375_));
 sky130_fd_sc_hd__nand2_1 _7046_ (.A(net368),
    .B(net2255),
    .Y(_3615_));
 sky130_fd_sc_hd__a21oi_1 _7047_ (.A1(_3607_),
    .A2(_3615_),
    .B1(net159),
    .Y(_1376_));
 sky130_fd_sc_hd__nand2_1 _7048_ (.A(net372),
    .B(_2700_),
    .Y(_3616_));
 sky130_fd_sc_hd__a21oi_1 _7049_ (.A1(_3607_),
    .A2(net2243),
    .B1(net159),
    .Y(_1377_));
 sky130_fd_sc_hd__nand2_1 _7050_ (.A(net386),
    .B(_2700_),
    .Y(_3617_));
 sky130_fd_sc_hd__a21oi_1 _7051_ (.A1(_3607_),
    .A2(net2239),
    .B1(net159),
    .Y(_1378_));
 sky130_fd_sc_hd__or2_1 _7052_ (.A(_1402_),
    .B(net1989),
    .X(_3618_));
 sky130_fd_sc_hd__a21oi_1 _7053_ (.A1(_3607_),
    .A2(_3618_),
    .B1(net159),
    .Y(_1379_));
 sky130_fd_sc_hd__nand2_1 _7054_ (.A(net694),
    .B(_2714_),
    .Y(_3619_));
 sky130_fd_sc_hd__or3b_4 _7055_ (.A(_2712_),
    .B(_2700_),
    .C_N(net2090),
    .X(_3620_));
 sky130_fd_sc_hd__a21oi_1 _7056_ (.A1(net695),
    .A2(_3620_),
    .B1(net159),
    .Y(_1380_));
 sky130_fd_sc_hd__nand2_1 _7057_ (.A(net399),
    .B(_2714_),
    .Y(_3621_));
 sky130_fd_sc_hd__a21oi_1 _7058_ (.A1(_3620_),
    .A2(_3621_),
    .B1(net159),
    .Y(_1381_));
 sky130_fd_sc_hd__nand2_1 _7059_ (.A(net402),
    .B(_2714_),
    .Y(_3622_));
 sky130_fd_sc_hd__a21oi_1 _7060_ (.A1(_3620_),
    .A2(_3622_),
    .B1(net159),
    .Y(_1382_));
 sky130_fd_sc_hd__nand2_1 _7061_ (.A(net409),
    .B(_2714_),
    .Y(_3623_));
 sky130_fd_sc_hd__a21oi_1 _7062_ (.A1(_3620_),
    .A2(_3623_),
    .B1(net159),
    .Y(_1383_));
 sky130_fd_sc_hd__nand2_1 _7063_ (.A(net419),
    .B(_2714_),
    .Y(_3624_));
 sky130_fd_sc_hd__a21oi_1 _7064_ (.A1(_3620_),
    .A2(_3624_),
    .B1(net159),
    .Y(_1384_));
 sky130_fd_sc_hd__nand2_1 _7065_ (.A(net2145),
    .B(_2714_),
    .Y(_3625_));
 sky130_fd_sc_hd__a21oi_1 _7066_ (.A1(_3620_),
    .A2(net2146),
    .B1(net160),
    .Y(_1385_));
 sky130_fd_sc_hd__nand2_1 _7067_ (.A(net1980),
    .B(_2714_),
    .Y(_3626_));
 sky130_fd_sc_hd__a21oi_1 _7068_ (.A1(_3620_),
    .A2(net1981),
    .B1(net160),
    .Y(_1386_));
 sky130_fd_sc_hd__nand2_1 _7069_ (.A(net2127),
    .B(_2714_),
    .Y(_3627_));
 sky130_fd_sc_hd__a21oi_1 _7070_ (.A1(_3620_),
    .A2(net2128),
    .B1(net160),
    .Y(_1387_));
 sky130_fd_sc_hd__nor2_1 _7071_ (.A(_2703_),
    .B(_3620_),
    .Y(_3628_));
 sky130_fd_sc_hd__a221o_1 _7072_ (.A1(net1957),
    .A2(_2703_),
    .B1(_2712_),
    .B2(net396),
    .C1(_3628_),
    .X(_3629_));
 sky130_fd_sc_hd__and3_1 _7073_ (.A(net179),
    .B(net232),
    .C(_3629_),
    .X(_1388_));
 sky130_fd_sc_hd__and3_1 _7074_ (.A(net2048),
    .B(_2679_),
    .C(net1989),
    .X(_1389_));
 sky130_fd_sc_hd__and3_1 _7075_ (.A(net1971),
    .B(_2679_),
    .C(net1989),
    .X(_1390_));
 sky130_fd_sc_hd__and3_1 _7076_ (.A(net2175),
    .B(_2679_),
    .C(net1989),
    .X(_1391_));
 sky130_fd_sc_hd__and3_1 _7077_ (.A(net1878),
    .B(_2679_),
    .C(net1989),
    .X(_1392_));
 sky130_fd_sc_hd__and3_1 _7078_ (.A(net2188),
    .B(_2679_),
    .C(net1989),
    .X(_1393_));
 sky130_fd_sc_hd__and3_1 _7079_ (.A(net2083),
    .B(_2679_),
    .C(net1989),
    .X(_1394_));
 sky130_fd_sc_hd__a21o_1 _7080_ (.A1(_2699_),
    .A2(net2171),
    .B1(_2712_),
    .X(_3630_));
 sky130_fd_sc_hd__a22o_1 _7081_ (.A1(net2198),
    .A2(_2701_),
    .B1(_3630_),
    .B2(net2109),
    .X(_3631_));
 sky130_fd_sc_hd__and3_1 _7082_ (.A(net176),
    .B(net225),
    .C(_3631_),
    .X(_1395_));
 sky130_fd_sc_hd__a22o_1 _7083_ (.A1(net2118),
    .A2(_2701_),
    .B1(_3630_),
    .B2(net2181),
    .X(_3632_));
 sky130_fd_sc_hd__and3_1 _7084_ (.A(net177),
    .B(net228),
    .C(net2182),
    .X(_1396_));
 sky130_fd_sc_hd__a22o_1 _7085_ (.A1(net2121),
    .A2(_2701_),
    .B1(_3630_),
    .B2(net375),
    .X(_3633_));
 sky130_fd_sc_hd__and3_1 _7086_ (.A(net177),
    .B(net228),
    .C(_3633_),
    .X(_1397_));
 sky130_fd_sc_hd__a22o_1 _7087_ (.A1(net1991),
    .A2(_2701_),
    .B1(_3630_),
    .B2(net386),
    .X(_3634_));
 sky130_fd_sc_hd__and3_1 _7088_ (.A(net177),
    .B(net228),
    .C(_3634_),
    .X(_1398_));
 sky130_fd_sc_hd__o32a_1 _7089_ (.A1(_1402_),
    .A2(_2701_),
    .A3(_2714_),
    .B1(_2711_),
    .B2(_1404_),
    .X(_3635_));
 sky130_fd_sc_hd__nor2_1 _7090_ (.A(net160),
    .B(net2172),
    .Y(_1399_));
 sky130_fd_sc_hd__o21a_1 _7091_ (.A1(_2174_),
    .A2(_2177_),
    .B1(_2176_),
    .X(_3637_));
 sky130_fd_sc_hd__o21a_1 _7092_ (.A1(_2174_),
    .A2(_2177_),
    .B1(_2176_),
    .X(_3638_));
 sky130_fd_sc_hd__o21a_1 _7093_ (.A1(_2174_),
    .A2(_2177_),
    .B1(_2176_),
    .X(_3639_));
 sky130_fd_sc_hd__o21a_1 _7094_ (.A1(_2174_),
    .A2(_2177_),
    .B1(_2176_),
    .X(_3640_));
 sky130_fd_sc_hd__inv_2 _7095_ (.A(net468),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _7096_ (.A(net464),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _7097_ (.A(net468),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _7098_ (.A(net468),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _7099_ (.A(net468),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _7100_ (.A(net468),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _7101_ (.A(net469),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _7102_ (.A(net468),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _7103_ (.A(net469),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _7104_ (.A(net469),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _7105_ (.A(net469),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _7106_ (.A(net469),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _7107_ (.A(net461),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _7108_ (.A(net461),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _7109_ (.A(net461),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _7110_ (.A(net463),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _7111_ (.A(net463),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _7112_ (.A(net463),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _7113_ (.A(net463),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _7114_ (.A(net461),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _7115_ (.A(net461),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _7116_ (.A(net463),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _7117_ (.A(net463),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _7118_ (.A(net465),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _7119_ (.A(net464),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _7120_ (.A(net464),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _7121_ (.A(net465),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _7122_ (.A(net464),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _7123_ (.A(net464),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _7124__2 (.A(clknet_leaf_50_clk),
    .Y(net478));
 sky130_fd_sc_hd__inv_2 _7125__3 (.A(clknet_leaf_43_clk),
    .Y(net479));
 sky130_fd_sc_hd__inv_2 _7126__4 (.A(clknet_leaf_42_clk),
    .Y(net480));
 sky130_fd_sc_hd__inv_2 _7127__5 (.A(clknet_leaf_95_clk),
    .Y(net481));
 sky130_fd_sc_hd__inv_2 _7128__6 (.A(clknet_leaf_25_clk),
    .Y(net482));
 sky130_fd_sc_hd__inv_2 _7129__7 (.A(clknet_leaf_26_clk),
    .Y(net483));
 sky130_fd_sc_hd__inv_2 _7130__8 (.A(clknet_leaf_101_clk),
    .Y(net484));
 sky130_fd_sc_hd__inv_2 _7131__9 (.A(clknet_leaf_49_clk),
    .Y(net485));
 sky130_fd_sc_hd__inv_2 _7132__10 (.A(clknet_leaf_26_clk),
    .Y(net486));
 sky130_fd_sc_hd__inv_2 _7133__11 (.A(clknet_leaf_33_clk),
    .Y(net487));
 sky130_fd_sc_hd__inv_2 _7134__12 (.A(clknet_leaf_9_clk),
    .Y(net488));
 sky130_fd_sc_hd__inv_2 _7135__13 (.A(clknet_leaf_35_clk),
    .Y(net489));
 sky130_fd_sc_hd__inv_2 _7136__14 (.A(clknet_leaf_43_clk),
    .Y(net490));
 sky130_fd_sc_hd__inv_2 _7137__15 (.A(clknet_leaf_18_clk),
    .Y(net491));
 sky130_fd_sc_hd__inv_2 _7138__16 (.A(clknet_leaf_2_clk),
    .Y(net492));
 sky130_fd_sc_hd__inv_2 _7139__17 (.A(clknet_leaf_7_clk),
    .Y(net493));
 sky130_fd_sc_hd__inv_2 _7140__18 (.A(clknet_leaf_42_clk),
    .Y(net494));
 sky130_fd_sc_hd__inv_2 _7141__19 (.A(clknet_leaf_2_clk),
    .Y(net495));
 sky130_fd_sc_hd__inv_2 _7142__20 (.A(clknet_leaf_7_clk),
    .Y(net496));
 sky130_fd_sc_hd__inv_2 _7143__21 (.A(clknet_leaf_1_clk),
    .Y(net497));
 sky130_fd_sc_hd__inv_2 _7144__22 (.A(clknet_leaf_20_clk),
    .Y(net498));
 sky130_fd_sc_hd__inv_2 _7145__23 (.A(clknet_leaf_103_clk),
    .Y(net499));
 sky130_fd_sc_hd__inv_2 _7146__24 (.A(clknet_leaf_112_clk),
    .Y(net500));
 sky130_fd_sc_hd__inv_2 _7147__25 (.A(clknet_leaf_96_clk),
    .Y(net501));
 sky130_fd_sc_hd__inv_2 _7148__26 (.A(clknet_leaf_8_clk),
    .Y(net502));
 sky130_fd_sc_hd__inv_2 _7149__27 (.A(clknet_leaf_111_clk),
    .Y(net503));
 sky130_fd_sc_hd__inv_2 _7150__28 (.A(clknet_leaf_105_clk),
    .Y(net504));
 sky130_fd_sc_hd__inv_2 _7151__29 (.A(clknet_leaf_11_clk),
    .Y(net505));
 sky130_fd_sc_hd__inv_2 _7152__30 (.A(clknet_leaf_100_clk),
    .Y(net506));
 sky130_fd_sc_hd__inv_2 _7153__31 (.A(clknet_leaf_10_clk),
    .Y(net507));
 sky130_fd_sc_hd__inv_2 _7154__32 (.A(clknet_leaf_14_clk),
    .Y(net508));
 sky130_fd_sc_hd__inv_2 _7155__33 (.A(clknet_leaf_86_clk),
    .Y(net509));
 sky130_fd_sc_hd__inv_2 _7156__34 (.A(clknet_leaf_4_clk),
    .Y(net510));
 sky130_fd_sc_hd__inv_2 _7157__35 (.A(clknet_leaf_94_clk),
    .Y(net511));
 sky130_fd_sc_hd__inv_2 _7158__36 (.A(clknet_leaf_6_clk),
    .Y(net512));
 sky130_fd_sc_hd__inv_2 _7159__37 (.A(clknet_leaf_54_clk),
    .Y(net513));
 sky130_fd_sc_hd__inv_2 _7160__38 (.A(clknet_leaf_30_clk),
    .Y(net514));
 sky130_fd_sc_hd__inv_2 _7161__39 (.A(clknet_leaf_32_clk),
    .Y(net515));
 sky130_fd_sc_hd__inv_2 _7162__40 (.A(clknet_leaf_92_clk),
    .Y(net516));
 sky130_fd_sc_hd__inv_2 _7163__41 (.A(clknet_leaf_23_clk),
    .Y(net517));
 sky130_fd_sc_hd__inv_2 _7164__42 (.A(clknet_leaf_29_clk),
    .Y(net518));
 sky130_fd_sc_hd__inv_2 _7165__43 (.A(clknet_leaf_59_clk),
    .Y(net519));
 sky130_fd_sc_hd__inv_2 _7166__44 (.A(clknet_leaf_28_clk),
    .Y(net520));
 sky130_fd_sc_hd__inv_2 _7167__45 (.A(clknet_leaf_28_clk),
    .Y(net521));
 sky130_fd_sc_hd__inv_2 _7168__46 (.A(clknet_leaf_0_clk),
    .Y(net522));
 sky130_fd_sc_hd__inv_2 _7169__47 (.A(clknet_leaf_115_clk),
    .Y(net523));
 sky130_fd_sc_hd__inv_2 _7170__48 (.A(clknet_leaf_115_clk),
    .Y(net524));
 sky130_fd_sc_hd__inv_2 _7171__49 (.A(clknet_leaf_5_clk),
    .Y(net525));
 sky130_fd_sc_hd__inv_2 _7172__50 (.A(clknet_leaf_36_clk),
    .Y(net526));
 sky130_fd_sc_hd__inv_2 _7173__51 (.A(clknet_leaf_52_clk),
    .Y(net527));
 sky130_fd_sc_hd__inv_2 _7174__52 (.A(clknet_leaf_6_clk),
    .Y(net528));
 sky130_fd_sc_hd__inv_2 _7175__53 (.A(clknet_leaf_115_clk),
    .Y(net529));
 sky130_fd_sc_hd__inv_2 _7176__54 (.A(clknet_leaf_0_clk),
    .Y(net530));
 sky130_fd_sc_hd__inv_2 _7177__55 (.A(clknet_leaf_52_clk),
    .Y(net531));
 sky130_fd_sc_hd__inv_2 _7178__56 (.A(clknet_leaf_94_clk),
    .Y(net532));
 sky130_fd_sc_hd__inv_2 _7179__57 (.A(clknet_leaf_59_clk),
    .Y(net533));
 sky130_fd_sc_hd__inv_2 _7180__58 (.A(clknet_leaf_85_clk),
    .Y(net534));
 sky130_fd_sc_hd__inv_2 _7181__59 (.A(clknet_leaf_115_clk),
    .Y(net535));
 sky130_fd_sc_hd__inv_2 _7182__60 (.A(clknet_leaf_115_clk),
    .Y(net536));
 sky130_fd_sc_hd__inv_2 _7183__61 (.A(clknet_leaf_114_clk),
    .Y(net537));
 sky130_fd_sc_hd__inv_2 _7184__62 (.A(clknet_leaf_108_clk),
    .Y(net538));
 sky130_fd_sc_hd__inv_2 _7185__63 (.A(clknet_leaf_66_clk),
    .Y(net539));
 sky130_fd_sc_hd__inv_2 _7186__64 (.A(clknet_leaf_94_clk),
    .Y(net540));
 sky130_fd_sc_hd__inv_2 _7187__65 (.A(clknet_leaf_115_clk),
    .Y(net541));
 sky130_fd_sc_hd__inv_2 _7188__66 (.A(clknet_leaf_56_clk),
    .Y(net542));
 sky130_fd_sc_hd__inv_2 _7189__67 (.A(clknet_leaf_47_clk),
    .Y(net543));
 sky130_fd_sc_hd__inv_2 _7190__68 (.A(clknet_leaf_43_clk),
    .Y(net544));
 sky130_fd_sc_hd__inv_2 _7191__69 (.A(clknet_leaf_43_clk),
    .Y(net545));
 sky130_fd_sc_hd__inv_2 _7192__70 (.A(clknet_leaf_82_clk),
    .Y(net546));
 sky130_fd_sc_hd__inv_2 _7193__71 (.A(clknet_leaf_17_clk),
    .Y(net547));
 sky130_fd_sc_hd__inv_2 _7194__72 (.A(clknet_leaf_34_clk),
    .Y(net548));
 sky130_fd_sc_hd__inv_2 _7195__73 (.A(clknet_leaf_70_clk),
    .Y(net549));
 sky130_fd_sc_hd__inv_2 _7196__74 (.A(clknet_leaf_63_clk),
    .Y(net550));
 sky130_fd_sc_hd__inv_2 _7197__75 (.A(clknet_leaf_47_clk),
    .Y(net551));
 sky130_fd_sc_hd__inv_2 _7198__76 (.A(clknet_leaf_50_clk),
    .Y(net552));
 sky130_fd_sc_hd__inv_2 _7199__77 (.A(clknet_leaf_12_clk),
    .Y(net553));
 sky130_fd_sc_hd__inv_2 _7200__78 (.A(clknet_leaf_55_clk),
    .Y(net554));
 sky130_fd_sc_hd__inv_2 _7201__79 (.A(clknet_leaf_48_clk),
    .Y(net555));
 sky130_fd_sc_hd__inv_2 _7202__80 (.A(clknet_leaf_16_clk),
    .Y(net556));
 sky130_fd_sc_hd__inv_2 _7203__81 (.A(clknet_leaf_10_clk),
    .Y(net557));
 sky130_fd_sc_hd__inv_2 _7204__82 (.A(clknet_leaf_15_clk),
    .Y(net558));
 sky130_fd_sc_hd__inv_2 _7205__83 (.A(clknet_leaf_63_clk),
    .Y(net559));
 sky130_fd_sc_hd__inv_2 _7206__84 (.A(clknet_leaf_100_clk),
    .Y(net560));
 sky130_fd_sc_hd__inv_2 _7207__85 (.A(clknet_leaf_8_clk),
    .Y(net561));
 sky130_fd_sc_hd__inv_2 _7208__86 (.A(clknet_leaf_110_clk),
    .Y(net562));
 sky130_fd_sc_hd__inv_2 _7209__87 (.A(clknet_leaf_15_clk),
    .Y(net563));
 sky130_fd_sc_hd__inv_2 _7210__88 (.A(clknet_leaf_74_clk),
    .Y(net564));
 sky130_fd_sc_hd__inv_2 _7211__89 (.A(clknet_leaf_92_clk),
    .Y(net565));
 sky130_fd_sc_hd__inv_2 _7212__90 (.A(clknet_leaf_89_clk),
    .Y(net566));
 sky130_fd_sc_hd__inv_2 _7213__91 (.A(clknet_leaf_13_clk),
    .Y(net567));
 sky130_fd_sc_hd__inv_2 _7214__92 (.A(clknet_leaf_81_clk),
    .Y(net568));
 sky130_fd_sc_hd__inv_2 _7215__93 (.A(clknet_leaf_83_clk),
    .Y(net569));
 sky130_fd_sc_hd__inv_2 _7216__94 (.A(clknet_leaf_76_clk),
    .Y(net570));
 sky130_fd_sc_hd__inv_2 _7217__95 (.A(clknet_leaf_80_clk),
    .Y(net571));
 sky130_fd_sc_hd__inv_2 _7218__96 (.A(clknet_leaf_13_clk),
    .Y(net572));
 sky130_fd_sc_hd__inv_2 _7219__97 (.A(clknet_leaf_73_clk),
    .Y(net573));
 sky130_fd_sc_hd__inv_2 _7220__98 (.A(clknet_leaf_50_clk),
    .Y(net574));
 sky130_fd_sc_hd__inv_2 _7221__99 (.A(clknet_leaf_50_clk),
    .Y(net575));
 sky130_fd_sc_hd__inv_2 _7222__100 (.A(clknet_leaf_43_clk),
    .Y(net576));
 sky130_fd_sc_hd__inv_2 _7223__101 (.A(clknet_leaf_42_clk),
    .Y(net577));
 sky130_fd_sc_hd__inv_2 _7224__102 (.A(clknet_leaf_96_clk),
    .Y(net578));
 sky130_fd_sc_hd__inv_2 _7225__103 (.A(clknet_leaf_25_clk),
    .Y(net579));
 sky130_fd_sc_hd__inv_2 _7226__104 (.A(clknet_leaf_27_clk),
    .Y(net580));
 sky130_fd_sc_hd__inv_2 _7227__105 (.A(clknet_leaf_101_clk),
    .Y(net581));
 sky130_fd_sc_hd__inv_2 _7228__106 (.A(clknet_leaf_49_clk),
    .Y(net582));
 sky130_fd_sc_hd__inv_2 _7229__107 (.A(clknet_leaf_26_clk),
    .Y(net583));
 sky130_fd_sc_hd__inv_2 _7230__108 (.A(clknet_leaf_33_clk),
    .Y(net584));
 sky130_fd_sc_hd__inv_2 _7231__109 (.A(clknet_leaf_9_clk),
    .Y(net585));
 sky130_fd_sc_hd__inv_2 _7232__110 (.A(clknet_leaf_34_clk),
    .Y(net586));
 sky130_fd_sc_hd__inv_2 _7233__111 (.A(clknet_leaf_43_clk),
    .Y(net587));
 sky130_fd_sc_hd__inv_2 _7234__112 (.A(clknet_leaf_18_clk),
    .Y(net588));
 sky130_fd_sc_hd__inv_2 _7235__113 (.A(clknet_leaf_3_clk),
    .Y(net589));
 sky130_fd_sc_hd__inv_2 _7236__114 (.A(clknet_leaf_20_clk),
    .Y(net590));
 sky130_fd_sc_hd__inv_2 _7237__115 (.A(clknet_leaf_17_clk),
    .Y(net591));
 sky130_fd_sc_hd__inv_2 _7238__116 (.A(clknet_leaf_2_clk),
    .Y(net592));
 sky130_fd_sc_hd__inv_2 _7239__117 (.A(clknet_leaf_7_clk),
    .Y(net593));
 sky130_fd_sc_hd__inv_2 _7240__118 (.A(clknet_leaf_1_clk),
    .Y(net594));
 sky130_fd_sc_hd__inv_2 _7241__119 (.A(clknet_leaf_18_clk),
    .Y(net595));
 sky130_fd_sc_hd__inv_2 _7242__120 (.A(clknet_leaf_103_clk),
    .Y(net596));
 sky130_fd_sc_hd__inv_2 _7243__121 (.A(clknet_leaf_112_clk),
    .Y(net597));
 sky130_fd_sc_hd__inv_2 _7244__122 (.A(clknet_leaf_96_clk),
    .Y(net598));
 sky130_fd_sc_hd__inv_2 _7245__123 (.A(clknet_leaf_12_clk),
    .Y(net599));
 sky130_fd_sc_hd__inv_2 _7246__124 (.A(clknet_leaf_104_clk),
    .Y(net600));
 sky130_fd_sc_hd__inv_2 _7247__125 (.A(clknet_leaf_106_clk),
    .Y(net601));
 sky130_fd_sc_hd__inv_2 _7248__126 (.A(clknet_leaf_11_clk),
    .Y(net602));
 sky130_fd_sc_hd__inv_2 _7249__127 (.A(clknet_leaf_100_clk),
    .Y(net603));
 sky130_fd_sc_hd__inv_2 _7250__128 (.A(clknet_leaf_10_clk),
    .Y(net604));
 sky130_fd_sc_hd__inv_2 _7251__129 (.A(clknet_leaf_14_clk),
    .Y(net605));
 sky130_fd_sc_hd__inv_2 _7252_ (.A(net468),
    .Y(_0260_));
 sky130_fd_sc_hd__inv_2 _7253_ (.A(net468),
    .Y(_0261_));
 sky130_fd_sc_hd__inv_2 _7254_ (.A(net464),
    .Y(_0262_));
 sky130_fd_sc_hd__inv_2 _7255_ (.A(net464),
    .Y(_0263_));
 sky130_fd_sc_hd__inv_2 _7256_ (.A(net468),
    .Y(_0264_));
 sky130_fd_sc_hd__inv_2 _7257_ (.A(net468),
    .Y(_0265_));
 sky130_fd_sc_hd__inv_2 _7258_ (.A(net468),
    .Y(_0266_));
 sky130_fd_sc_hd__inv_2 _7259_ (.A(net469),
    .Y(_0267_));
 sky130_fd_sc_hd__inv_2 _7260_ (.A(net469),
    .Y(_0268_));
 sky130_fd_sc_hd__inv_2 _7261_ (.A(net469),
    .Y(_0269_));
 sky130_fd_sc_hd__inv_2 _7262_ (.A(net469),
    .Y(_0270_));
 sky130_fd_sc_hd__inv_2 _7263_ (.A(net469),
    .Y(_0271_));
 sky130_fd_sc_hd__inv_2 _7264_ (.A(net469),
    .Y(_0272_));
 sky130_fd_sc_hd__inv_2 _7265_ (.A(net461),
    .Y(_0273_));
 sky130_fd_sc_hd__inv_2 _7266_ (.A(net461),
    .Y(_0274_));
 sky130_fd_sc_hd__inv_2 _7267_ (.A(net461),
    .Y(_0275_));
 sky130_fd_sc_hd__inv_2 _7268_ (.A(net463),
    .Y(_0276_));
 sky130_fd_sc_hd__inv_2 _7269_ (.A(net463),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_2 _7270_ (.A(net463),
    .Y(_0278_));
 sky130_fd_sc_hd__inv_2 _7271_ (.A(net463),
    .Y(_0279_));
 sky130_fd_sc_hd__inv_2 _7272_ (.A(net463),
    .Y(_0280_));
 sky130_fd_sc_hd__inv_2 _7273_ (.A(net463),
    .Y(_0281_));
 sky130_fd_sc_hd__inv_2 _7274_ (.A(net465),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_2 _7275_ (.A(net465),
    .Y(_0283_));
 sky130_fd_sc_hd__inv_2 _7276_ (.A(net465),
    .Y(_0284_));
 sky130_fd_sc_hd__inv_2 _7277_ (.A(net464),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_2 _7278_ (.A(net464),
    .Y(_0286_));
 sky130_fd_sc_hd__inv_2 _7279_ (.A(net464),
    .Y(_0287_));
 sky130_fd_sc_hd__inv_2 _7280_ (.A(net465),
    .Y(_0288_));
 sky130_fd_sc_hd__inv_2 _7281_ (.A(net465),
    .Y(_0289_));
 sky130_fd_sc_hd__dfxtp_2 _7282_ (.CLK(clknet_leaf_56_clk),
    .D(net802),
    .Q(\U_DATAPATH.U_MEM_WB.o_result_src_WB[0] ));
 sky130_fd_sc_hd__dfxtp_4 _7283_ (.CLK(clknet_leaf_56_clk),
    .D(net744),
    .Q(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7284_ (.CLK(clknet_leaf_69_clk),
    .D(_0292_),
    .RESET_B(net452),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_1 _7285_ (.CLK(clknet_leaf_67_clk),
    .D(_0293_),
    .RESET_B(_0102_),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_4 _7286_ (.CLK(clknet_leaf_77_clk),
    .D(_0294_),
    .RESET_B(_0103_),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_4 _7287_ (.CLK(clknet_leaf_68_clk),
    .D(_0295_),
    .RESET_B(_0104_),
    .Q(net122));
 sky130_fd_sc_hd__dfrtp_2 _7288_ (.CLK(clknet_leaf_67_clk),
    .D(_0296_),
    .RESET_B(_0105_),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_4 _7289_ (.CLK(clknet_leaf_71_clk),
    .D(_0297_),
    .RESET_B(_0106_),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_1 _7290_ (.CLK(clknet_leaf_66_clk),
    .D(_0298_),
    .RESET_B(_0107_),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_2 _7291_ (.CLK(clknet_leaf_61_clk),
    .D(_0299_),
    .RESET_B(_0108_),
    .Q(net126));
 sky130_fd_sc_hd__dfrtp_4 _7292_ (.CLK(clknet_leaf_63_clk),
    .D(_0300_),
    .RESET_B(_0109_),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_4 _7293_ (.CLK(clknet_leaf_56_clk),
    .D(_0301_),
    .RESET_B(_0110_),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_4 _7294_ (.CLK(clknet_leaf_57_clk),
    .D(_0302_),
    .RESET_B(_0111_),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_4 _7295_ (.CLK(clknet_leaf_61_clk),
    .D(_0303_),
    .RESET_B(_0112_),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_2 _7296_ (.CLK(clknet_leaf_57_clk),
    .D(_0304_),
    .RESET_B(_0113_),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_4 _7297_ (.CLK(clknet_leaf_94_clk),
    .D(_0305_),
    .RESET_B(_0114_),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_4 _7298_ (.CLK(clknet_leaf_95_clk),
    .D(_0306_),
    .RESET_B(_0115_),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_4 _7299_ (.CLK(clknet_leaf_97_clk),
    .D(_0307_),
    .RESET_B(_0116_),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_4 _7300_ (.CLK(clknet_leaf_74_clk),
    .D(_0308_),
    .RESET_B(_0117_),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_2 _7301_ (.CLK(clknet_leaf_74_clk),
    .D(_0309_),
    .RESET_B(_0118_),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_4 _7302_ (.CLK(clknet_leaf_90_clk),
    .D(_0310_),
    .RESET_B(_0119_),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_4 _7303_ (.CLK(clknet_leaf_82_clk),
    .D(_0311_),
    .RESET_B(_0120_),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_4 _7304_ (.CLK(clknet_leaf_90_clk),
    .D(_0312_),
    .RESET_B(_0121_),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_4 _7305_ (.CLK(clknet_leaf_91_clk),
    .D(_0313_),
    .RESET_B(_0122_),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_1 _7306_ (.CLK(clknet_leaf_83_clk),
    .D(_0314_),
    .RESET_B(_0123_),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_2 _7307_ (.CLK(clknet_leaf_89_clk),
    .D(_0315_),
    .RESET_B(_0124_),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_2 _7308_ (.CLK(clknet_leaf_83_clk),
    .D(_0316_),
    .RESET_B(_0125_),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_4 _7309_ (.CLK(clknet_leaf_81_clk),
    .D(_0317_),
    .RESET_B(_0126_),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_2 _7310_ (.CLK(clknet_leaf_81_clk),
    .D(_0318_),
    .RESET_B(_0127_),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_4 _7311_ (.CLK(clknet_leaf_81_clk),
    .D(_0319_),
    .RESET_B(_0128_),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_4 _7312_ (.CLK(clknet_leaf_79_clk),
    .D(_0320_),
    .RESET_B(_0129_),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_4 _7313_ (.CLK(clknet_leaf_78_clk),
    .D(_0321_),
    .RESET_B(_0130_),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_1 _7314_ (.CLK(clknet_leaf_64_clk),
    .D(_0322_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7315_ (.CLK(clknet_leaf_68_clk),
    .D(_0323_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7316_ (.CLK(clknet_leaf_78_clk),
    .D(_0324_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7317_ (.CLK(clknet_leaf_78_clk),
    .D(net838),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7318_ (.CLK(clknet_leaf_66_clk),
    .D(net818),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7319_ (.CLK(clknet_leaf_69_clk),
    .D(_0327_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7320_ (.CLK(clknet_leaf_65_clk),
    .D(net1894),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7321_ (.CLK(clknet_leaf_65_clk),
    .D(_0329_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7322_ (.CLK(clknet_leaf_62_clk),
    .D(_0330_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7323_ (.CLK(clknet_leaf_57_clk),
    .D(_0331_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7324_ (.CLK(clknet_leaf_57_clk),
    .D(_0332_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7325_ (.CLK(clknet_leaf_60_clk),
    .D(net1793),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7326_ (.CLK(clknet_leaf_60_clk),
    .D(net1243),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7327_ (.CLK(clknet_leaf_93_clk),
    .D(_0335_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7328_ (.CLK(clknet_leaf_93_clk),
    .D(_0336_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7329_ (.CLK(clknet_leaf_91_clk),
    .D(_0337_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7330_ (.CLK(clknet_leaf_82_clk),
    .D(_0338_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7331_ (.CLK(clknet_leaf_98_clk),
    .D(net1785),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7332_ (.CLK(clknet_leaf_89_clk),
    .D(_0340_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7333_ (.CLK(clknet_leaf_98_clk),
    .D(_0341_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7334_ (.CLK(clknet_leaf_91_clk),
    .D(net1821),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7335_ (.CLK(clknet_leaf_91_clk),
    .D(_0343_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7336_ (.CLK(clknet_leaf_89_clk),
    .D(_0344_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7337_ (.CLK(clknet_leaf_83_clk),
    .D(_0345_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7338_ (.CLK(clknet_leaf_84_clk),
    .D(_0346_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7339_ (.CLK(clknet_leaf_79_clk),
    .D(net872),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7340_ (.CLK(clknet_leaf_75_clk),
    .D(_0348_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7341_ (.CLK(clknet_leaf_81_clk),
    .D(_0349_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7342_ (.CLK(clknet_leaf_79_clk),
    .D(_0350_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7343_ (.CLK(clknet_leaf_76_clk),
    .D(_0351_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7344_ (.CLK(clknet_leaf_59_clk),
    .D(_0352_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7345_ (.CLK(clknet_leaf_86_clk),
    .D(_0353_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7346_ (.CLK(clknet_leaf_88_clk),
    .D(_0354_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7347_ (.CLK(clknet_leaf_74_clk),
    .D(_0355_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7348_ (.CLK(clknet_leaf_66_clk),
    .D(_0356_),
    .Q(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7349_ (.CLK(clknet_leaf_47_clk),
    .D(_0357_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7350_ (.CLK(clknet_leaf_36_clk),
    .D(_0358_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7351_ (.CLK(clknet_leaf_53_clk),
    .D(_0359_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7352_ (.CLK(clknet_leaf_54_clk),
    .D(_0360_),
    .Q(\U_DATAPATH.U_ID_EX.i_rd_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7353_ (.CLK(clknet_leaf_66_clk),
    .D(_0361_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7354_ (.CLK(clknet_leaf_54_clk),
    .D(_0362_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7355_ (.CLK(clknet_leaf_73_clk),
    .D(_0363_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7356_ (.CLK(clknet_leaf_59_clk),
    .D(_0364_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ));
 sky130_fd_sc_hd__dfxtp_4 _7357_ (.CLK(clknet_leaf_114_clk),
    .D(_0365_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7358_ (.CLK(clknet_leaf_87_clk),
    .D(_0366_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7359_ (.CLK(clknet_leaf_53_clk),
    .D(_0367_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7360_ (.CLK(clknet_leaf_80_clk),
    .D(_0368_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7361_ (.CLK(clknet_leaf_68_clk),
    .D(_0369_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[19] ));
 sky130_fd_sc_hd__dfxtp_4 _7362_ (.CLK(clknet_leaf_9_clk),
    .D(_0370_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7363_ (.CLK(clknet_leaf_38_clk),
    .D(_0371_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7364_ (.CLK(clknet_leaf_114_clk),
    .D(_0372_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ));
 sky130_fd_sc_hd__dfxtp_4 _7365_ (.CLK(clknet_leaf_25_clk),
    .D(_0373_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7366_ (.CLK(clknet_leaf_94_clk),
    .D(_0374_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7367_ (.CLK(clknet_leaf_78_clk),
    .D(_0375_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7368_ (.CLK(clknet_leaf_31_clk),
    .D(_0376_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7369_ (.CLK(clknet_leaf_58_clk),
    .D(_0377_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7370_ (.CLK(clknet_leaf_18_clk),
    .D(_0378_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7371_ (.CLK(clknet_leaf_85_clk),
    .D(_0379_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7372_ (.CLK(clknet_leaf_56_clk),
    .D(_0380_),
    .Q(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ));
 sky130_fd_sc_hd__dfxtp_1 _7373_ (.CLK(clknet_leaf_54_clk),
    .D(_0381_),
    .Q(\U_DATAPATH.U_IF_ID.o_instr_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7374_ (.CLK(clknet_leaf_69_clk),
    .D(_0382_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7375_ (.CLK(clknet_leaf_67_clk),
    .D(_0383_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7376_ (.CLK(clknet_leaf_78_clk),
    .D(_0384_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7377_ (.CLK(clknet_leaf_70_clk),
    .D(_0385_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7378_ (.CLK(clknet_leaf_67_clk),
    .D(_0386_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7379_ (.CLK(clknet_leaf_71_clk),
    .D(_0387_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7380_ (.CLK(clknet_leaf_66_clk),
    .D(_0388_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7381_ (.CLK(clknet_leaf_61_clk),
    .D(_0389_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7382_ (.CLK(clknet_leaf_63_clk),
    .D(_0390_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7383_ (.CLK(clknet_leaf_56_clk),
    .D(_0391_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7384_ (.CLK(clknet_leaf_57_clk),
    .D(_0392_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7385_ (.CLK(clknet_leaf_61_clk),
    .D(_0393_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7386_ (.CLK(clknet_leaf_57_clk),
    .D(_0394_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7387_ (.CLK(clknet_leaf_95_clk),
    .D(_0395_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7388_ (.CLK(clknet_leaf_96_clk),
    .D(_0396_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7389_ (.CLK(clknet_leaf_98_clk),
    .D(_0397_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7390_ (.CLK(clknet_leaf_98_clk),
    .D(_0398_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7391_ (.CLK(clknet_leaf_82_clk),
    .D(_0399_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7392_ (.CLK(clknet_leaf_90_clk),
    .D(_0400_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7393_ (.CLK(clknet_leaf_82_clk),
    .D(_0401_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7394_ (.CLK(clknet_leaf_97_clk),
    .D(_0402_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7395_ (.CLK(clknet_leaf_91_clk),
    .D(_0403_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7396_ (.CLK(clknet_leaf_83_clk),
    .D(_0404_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7397_ (.CLK(clknet_leaf_89_clk),
    .D(_0405_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7398_ (.CLK(clknet_leaf_85_clk),
    .D(_0406_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7399_ (.CLK(clknet_leaf_74_clk),
    .D(_0407_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7400_ (.CLK(clknet_leaf_81_clk),
    .D(_0408_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7401_ (.CLK(clknet_leaf_74_clk),
    .D(_0409_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7402_ (.CLK(clknet_leaf_79_clk),
    .D(_0410_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7403_ (.CLK(clknet_leaf_78_clk),
    .D(_0411_),
    .Q(\U_DATAPATH.U_ID_EX.i_pc_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7404_ (.CLK(clknet_leaf_41_clk),
    .D(net1149),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7405_ (.CLK(clknet_leaf_41_clk),
    .D(net950),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7406_ (.CLK(clknet_leaf_35_clk),
    .D(net892),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7407_ (.CLK(clknet_leaf_35_clk),
    .D(net890),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7408_ (.CLK(clknet_leaf_106_clk),
    .D(net1689),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7409_ (.CLK(clknet_leaf_23_clk),
    .D(net1079),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7410_ (.CLK(clknet_leaf_27_clk),
    .D(net1273),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7411_ (.CLK(clknet_leaf_11_clk),
    .D(net1639),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7412_ (.CLK(clknet_leaf_43_clk),
    .D(net1647),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7413_ (.CLK(clknet_leaf_27_clk),
    .D(net1427),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7414_ (.CLK(clknet_leaf_26_clk),
    .D(net1463),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7415_ (.CLK(clknet_leaf_5_clk),
    .D(net1227),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7416_ (.CLK(clknet_leaf_34_clk),
    .D(net1275),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7417_ (.CLK(clknet_leaf_17_clk),
    .D(net1537),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7418_ (.CLK(clknet_leaf_18_clk),
    .D(net1357),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7419_ (.CLK(clknet_leaf_4_clk),
    .D(net1111),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7420_ (.CLK(clknet_leaf_21_clk),
    .D(net1053),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7421_ (.CLK(clknet_leaf_26_clk),
    .D(net1415),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7422_ (.CLK(clknet_leaf_1_clk),
    .D(net1439),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7423_ (.CLK(clknet_leaf_7_clk),
    .D(net1603),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7424_ (.CLK(clknet_leaf_0_clk),
    .D(net1279),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7425_ (.CLK(clknet_leaf_23_clk),
    .D(net1245),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7426_ (.CLK(clknet_leaf_10_clk),
    .D(net1455),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7427_ (.CLK(clknet_leaf_112_clk),
    .D(net1215),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7428_ (.CLK(clknet_leaf_105_clk),
    .D(net1209),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7429_ (.CLK(clknet_leaf_20_clk),
    .D(net1365),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7430_ (.CLK(clknet_leaf_112_clk),
    .D(net1107),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7431_ (.CLK(clknet_leaf_105_clk),
    .D(net1073),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7432_ (.CLK(clknet_leaf_11_clk),
    .D(net1561),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7433_ (.CLK(clknet_leaf_102_clk),
    .D(net1623),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7434_ (.CLK(clknet_leaf_9_clk),
    .D(net1341),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7435_ (.CLK(clknet_leaf_14_clk),
    .D(net1523),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7436_ (.CLK(clknet_leaf_37_clk),
    .D(net940),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7437_ (.CLK(clknet_leaf_37_clk),
    .D(net964),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7438_ (.CLK(clknet_leaf_42_clk),
    .D(net1381),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7439_ (.CLK(clknet_leaf_37_clk),
    .D(net860),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7440_ (.CLK(clknet_leaf_107_clk),
    .D(net1465),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7441_ (.CLK(clknet_leaf_25_clk),
    .D(net1359),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7442_ (.CLK(clknet_leaf_29_clk),
    .D(net1407),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7443_ (.CLK(clknet_leaf_103_clk),
    .D(net1595),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7444_ (.CLK(clknet_leaf_41_clk),
    .D(net1479),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7445_ (.CLK(clknet_leaf_27_clk),
    .D(net1151),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7446_ (.CLK(clknet_leaf_33_clk),
    .D(net1123),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7447_ (.CLK(clknet_leaf_3_clk),
    .D(net1255),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7448_ (.CLK(clknet_leaf_33_clk),
    .D(net1201),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7449_ (.CLK(clknet_leaf_42_clk),
    .D(net1713),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7450_ (.CLK(clknet_leaf_18_clk),
    .D(net1095),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7451_ (.CLK(clknet_leaf_0_clk),
    .D(net1213),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7452_ (.CLK(clknet_leaf_6_clk),
    .D(net1025),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7453_ (.CLK(clknet_leaf_26_clk),
    .D(net1533),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7454_ (.CLK(clknet_leaf_1_clk),
    .D(net1087),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7455_ (.CLK(clknet_leaf_7_clk),
    .D(net1581),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7456_ (.CLK(clknet_leaf_116_clk),
    .D(net1000),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7457_ (.CLK(clknet_leaf_21_clk),
    .D(net1035),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7458_ (.CLK(clknet_leaf_10_clk),
    .D(net1283),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7459_ (.CLK(clknet_leaf_113_clk),
    .D(net1141),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7460_ (.CLK(clknet_leaf_105_clk),
    .D(net1055),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7461_ (.CLK(clknet_leaf_19_clk),
    .D(net982),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7462_ (.CLK(clknet_leaf_111_clk),
    .D(net1155),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7463_ (.CLK(clknet_leaf_111_clk),
    .D(net1059),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7464_ (.CLK(clknet_leaf_11_clk),
    .D(net1307),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7465_ (.CLK(clknet_leaf_106_clk),
    .D(net1651),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7466_ (.CLK(clknet_leaf_3_clk),
    .D(net1085),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7467_ (.CLK(clknet_leaf_15_clk),
    .D(net1573),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7468_ (.CLK(clknet_leaf_39_clk),
    .D(net958),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7469_ (.CLK(clknet_leaf_39_clk),
    .D(net906),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7470_ (.CLK(clknet_leaf_42_clk),
    .D(net1667),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7471_ (.CLK(clknet_leaf_39_clk),
    .D(net836),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7472_ (.CLK(clknet_leaf_107_clk),
    .D(net1655),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7473_ (.CLK(clknet_leaf_24_clk),
    .D(net1147),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7474_ (.CLK(clknet_leaf_29_clk),
    .D(net1393),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7475_ (.CLK(clknet_leaf_103_clk),
    .D(net1699),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7476_ (.CLK(clknet_leaf_41_clk),
    .D(net1387),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7477_ (.CLK(clknet_leaf_25_clk),
    .D(net1571),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7478_ (.CLK(clknet_leaf_33_clk),
    .D(net1203),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7479_ (.CLK(clknet_leaf_3_clk),
    .D(net1429),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7480_ (.CLK(clknet_leaf_33_clk),
    .D(net1271),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7481_ (.CLK(clknet_leaf_42_clk),
    .D(net1585),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7482_ (.CLK(clknet_leaf_20_clk),
    .D(net1529),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7483_ (.CLK(clknet_leaf_0_clk),
    .D(net1235),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7484_ (.CLK(clknet_leaf_6_clk),
    .D(net1129),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7485_ (.CLK(clknet_leaf_25_clk),
    .D(net1643),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7486_ (.CLK(clknet_leaf_113_clk),
    .D(net1183),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7487_ (.CLK(clknet_leaf_5_clk),
    .D(net1247),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7488_ (.CLK(clknet_leaf_116_clk),
    .D(net1127),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7489_ (.CLK(clknet_leaf_21_clk),
    .D(net1417),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7490_ (.CLK(clknet_leaf_10_clk),
    .D(net1397),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7491_ (.CLK(clknet_leaf_113_clk),
    .D(net1421),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7492_ (.CLK(clknet_leaf_105_clk),
    .D(net1285),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7493_ (.CLK(clknet_leaf_19_clk),
    .D(net978),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7494_ (.CLK(clknet_leaf_111_clk),
    .D(net1169),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7495_ (.CLK(clknet_leaf_111_clk),
    .D(net1351),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7496_ (.CLK(clknet_leaf_11_clk),
    .D(net1353),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7497_ (.CLK(clknet_leaf_106_clk),
    .D(net1663),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7498_ (.CLK(clknet_leaf_3_clk),
    .D(net1125),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7499_ (.CLK(clknet_leaf_15_clk),
    .D(net1467),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7500_ (.CLK(net477),
    .D(_0000_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7501_ (.CLK(net478),
    .D(_0011_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7502_ (.CLK(net479),
    .D(_0022_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7503_ (.CLK(net480),
    .D(_0025_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7504_ (.CLK(net481),
    .D(_0026_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7505_ (.CLK(net482),
    .D(_0027_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7506_ (.CLK(net483),
    .D(_0028_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7507_ (.CLK(net484),
    .D(_0029_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7508_ (.CLK(net485),
    .D(_0030_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7509_ (.CLK(net486),
    .D(_0031_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7510_ (.CLK(net487),
    .D(_0001_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7511_ (.CLK(net488),
    .D(_0002_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7512_ (.CLK(net489),
    .D(_0003_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7513_ (.CLK(net490),
    .D(_0004_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7514_ (.CLK(net491),
    .D(_0005_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7515_ (.CLK(net492),
    .D(_0006_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7516_ (.CLK(net493),
    .D(_0007_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7517_ (.CLK(net494),
    .D(_0008_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7518_ (.CLK(net495),
    .D(_0009_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7519_ (.CLK(net496),
    .D(_0010_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7520_ (.CLK(net497),
    .D(_0012_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7521_ (.CLK(net498),
    .D(_0013_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7522_ (.CLK(net499),
    .D(_0014_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7523_ (.CLK(net500),
    .D(_0015_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7524_ (.CLK(net501),
    .D(_0016_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7525_ (.CLK(net502),
    .D(_0017_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7526_ (.CLK(net503),
    .D(_0018_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7527_ (.CLK(net504),
    .D(_0019_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7528_ (.CLK(net505),
    .D(_0020_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7529_ (.CLK(net506),
    .D(_0021_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7530_ (.CLK(net507),
    .D(_0023_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7531_ (.CLK(net508),
    .D(_0024_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs2_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7532_ (.CLK(clknet_leaf_41_clk),
    .D(net870),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7533_ (.CLK(clknet_leaf_40_clk),
    .D(net1069),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7534_ (.CLK(clknet_leaf_41_clk),
    .D(net844),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7535_ (.CLK(clknet_leaf_41_clk),
    .D(net966),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7536_ (.CLK(clknet_leaf_106_clk),
    .D(net1331),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7537_ (.CLK(clknet_leaf_25_clk),
    .D(net1389),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7538_ (.CLK(clknet_leaf_27_clk),
    .D(net1471),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7539_ (.CLK(clknet_leaf_13_clk),
    .D(net1773),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7540_ (.CLK(clknet_leaf_44_clk),
    .D(net1027),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7541_ (.CLK(clknet_leaf_26_clk),
    .D(net1635),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7542_ (.CLK(clknet_leaf_34_clk),
    .D(net1019),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7543_ (.CLK(clknet_leaf_3_clk),
    .D(net1004),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7544_ (.CLK(clknet_leaf_35_clk),
    .D(net1683),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7545_ (.CLK(clknet_leaf_42_clk),
    .D(net1521),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7546_ (.CLK(clknet_leaf_17_clk),
    .D(net1513),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7547_ (.CLK(clknet_leaf_3_clk),
    .D(net1117),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7548_ (.CLK(clknet_leaf_20_clk),
    .D(net1199),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7549_ (.CLK(clknet_leaf_42_clk),
    .D(net1601),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7550_ (.CLK(clknet_leaf_1_clk),
    .D(net1233),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7551_ (.CLK(clknet_leaf_7_clk),
    .D(net1563),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7552_ (.CLK(clknet_leaf_0_clk),
    .D(net1691),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7553_ (.CLK(clknet_leaf_18_clk),
    .D(net1077),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7554_ (.CLK(clknet_leaf_11_clk),
    .D(net1299),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7555_ (.CLK(clknet_leaf_112_clk),
    .D(net1507),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7556_ (.CLK(clknet_leaf_105_clk),
    .D(net1319),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7557_ (.CLK(clknet_leaf_20_clk),
    .D(net1383),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7558_ (.CLK(clknet_leaf_104_clk),
    .D(net1555),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7559_ (.CLK(clknet_leaf_104_clk),
    .D(net1503),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7560_ (.CLK(clknet_leaf_13_clk),
    .D(net1591),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7561_ (.CLK(clknet_leaf_102_clk),
    .D(net1016),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7562_ (.CLK(clknet_leaf_9_clk),
    .D(net1137),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7563_ (.CLK(clknet_leaf_14_clk),
    .D(net1093),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7564_ (.CLK(clknet_leaf_39_clk),
    .D(net834),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7565_ (.CLK(clknet_leaf_39_clk),
    .D(net852),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7566_ (.CLK(clknet_leaf_41_clk),
    .D(net864),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7567_ (.CLK(clknet_leaf_35_clk),
    .D(net896),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7568_ (.CLK(clknet_leaf_105_clk),
    .D(net1661),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7569_ (.CLK(clknet_leaf_25_clk),
    .D(net1525),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7570_ (.CLK(clknet_leaf_27_clk),
    .D(net1229),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7571_ (.CLK(clknet_leaf_11_clk),
    .D(net1565),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7572_ (.CLK(clknet_leaf_43_clk),
    .D(net1645),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7573_ (.CLK(clknet_leaf_27_clk),
    .D(net1021),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7574_ (.CLK(clknet_leaf_26_clk),
    .D(net1505),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7575_ (.CLK(clknet_leaf_5_clk),
    .D(net1163),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7576_ (.CLK(clknet_leaf_34_clk),
    .D(net1631),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7577_ (.CLK(clknet_leaf_17_clk),
    .D(net1583),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7578_ (.CLK(clknet_leaf_18_clk),
    .D(net1481),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7579_ (.CLK(clknet_leaf_4_clk),
    .D(net1167),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7580_ (.CLK(clknet_leaf_21_clk),
    .D(net1008),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7581_ (.CLK(clknet_leaf_26_clk),
    .D(net1413),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7582_ (.CLK(clknet_leaf_1_clk),
    .D(net1173),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7583_ (.CLK(clknet_leaf_7_clk),
    .D(net1305),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7584_ (.CLK(clknet_leaf_0_clk),
    .D(net1355),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7585_ (.CLK(clknet_leaf_23_clk),
    .D(net1047),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7586_ (.CLK(clknet_leaf_10_clk),
    .D(net1551),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7587_ (.CLK(clknet_leaf_112_clk),
    .D(net1121),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7588_ (.CLK(clknet_leaf_105_clk),
    .D(net1029),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7589_ (.CLK(clknet_leaf_20_clk),
    .D(net1221),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7590_ (.CLK(clknet_leaf_112_clk),
    .D(net1165),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7591_ (.CLK(clknet_leaf_104_clk),
    .D(net1419),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7592_ (.CLK(clknet_leaf_11_clk),
    .D(net1395),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7593_ (.CLK(clknet_leaf_102_clk),
    .D(net1375),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7594_ (.CLK(clknet_leaf_3_clk),
    .D(net1159),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7595_ (.CLK(clknet_leaf_14_clk),
    .D(net1317),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7596_ (.CLK(clknet_leaf_70_clk),
    .D(_0572_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7597_ (.CLK(clknet_leaf_92_clk),
    .D(_0573_),
    .Q(\U_DATAPATH.U_EX_MEM.i_mem_write_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7598_ (.CLK(clknet_leaf_56_clk),
    .D(_0574_),
    .Q(\U_DATAPATH.U_EX_MEM.i_result_src_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7599_ (.CLK(clknet_leaf_56_clk),
    .D(_0575_),
    .Q(\U_DATAPATH.U_EX_MEM.i_reg_write_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7600_ (.CLK(clknet_leaf_64_clk),
    .D(net926),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7601_ (.CLK(clknet_leaf_68_clk),
    .D(net1014),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7602_ (.CLK(clknet_leaf_77_clk),
    .D(net840),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7603_ (.CLK(clknet_leaf_78_clk),
    .D(net936),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7604_ (.CLK(clknet_leaf_66_clk),
    .D(net920),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7605_ (.CLK(clknet_leaf_69_clk),
    .D(net884),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7606_ (.CLK(clknet_leaf_65_clk),
    .D(net898),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7607_ (.CLK(clknet_leaf_65_clk),
    .D(net970),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7608_ (.CLK(clknet_leaf_62_clk),
    .D(net878),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7609_ (.CLK(clknet_leaf_54_clk),
    .D(net850),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7610_ (.CLK(clknet_leaf_57_clk),
    .D(net932),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7611_ (.CLK(clknet_leaf_60_clk),
    .D(net944),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7612_ (.CLK(clknet_leaf_60_clk),
    .D(net974),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7613_ (.CLK(clknet_leaf_93_clk),
    .D(net1153),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7614_ (.CLK(clknet_leaf_93_clk),
    .D(net922),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7615_ (.CLK(clknet_leaf_91_clk),
    .D(net952),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7616_ (.CLK(clknet_leaf_82_clk),
    .D(net986),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7617_ (.CLK(clknet_leaf_98_clk),
    .D(net1323),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7618_ (.CLK(clknet_leaf_88_clk),
    .D(net810),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7619_ (.CLK(clknet_leaf_97_clk),
    .D(net784),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7620_ (.CLK(clknet_leaf_92_clk),
    .D(net804),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7621_ (.CLK(clknet_leaf_92_clk),
    .D(net822),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7622_ (.CLK(clknet_leaf_87_clk),
    .D(net902),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7623_ (.CLK(clknet_leaf_81_clk),
    .D(net704),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7624_ (.CLK(clknet_leaf_84_clk),
    .D(net894),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7625_ (.CLK(clknet_leaf_79_clk),
    .D(net946),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7626_ (.CLK(clknet_leaf_75_clk),
    .D(net914),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7627_ (.CLK(clknet_leaf_81_clk),
    .D(net956),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7628_ (.CLK(clknet_leaf_79_clk),
    .D(net990),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7629_ (.CLK(clknet_leaf_76_clk),
    .D(net942),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7630_ (.CLK(clknet_leaf_69_clk),
    .D(net888),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7631_ (.CLK(clknet_leaf_67_clk),
    .D(net874),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7632_ (.CLK(clknet_leaf_77_clk),
    .D(net820),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7633_ (.CLK(clknet_leaf_69_clk),
    .D(net828),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7634_ (.CLK(clknet_leaf_67_clk),
    .D(net1131),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7635_ (.CLK(clknet_leaf_71_clk),
    .D(net876),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7636_ (.CLK(clknet_leaf_64_clk),
    .D(net854),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7637_ (.CLK(clknet_leaf_65_clk),
    .D(net824),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7638_ (.CLK(clknet_leaf_63_clk),
    .D(net962),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7639_ (.CLK(clknet_leaf_56_clk),
    .D(net988),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7640_ (.CLK(clknet_leaf_57_clk),
    .D(net938),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7641_ (.CLK(clknet_leaf_61_clk),
    .D(net900),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7642_ (.CLK(clknet_leaf_62_clk),
    .D(net968),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7643_ (.CLK(clknet_leaf_97_clk),
    .D(net996),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7644_ (.CLK(clknet_leaf_96_clk),
    .D(net980),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7645_ (.CLK(clknet_leaf_98_clk),
    .D(net994),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7646_ (.CLK(clknet_leaf_74_clk),
    .D(net814),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7647_ (.CLK(clknet_leaf_82_clk),
    .D(net1105),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7648_ (.CLK(clknet_leaf_90_clk),
    .D(net916),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7649_ (.CLK(clknet_leaf_89_clk),
    .D(net649),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7650_ (.CLK(clknet_leaf_97_clk),
    .D(net856),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7651_ (.CLK(clknet_leaf_91_clk),
    .D(net930),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7652_ (.CLK(clknet_leaf_83_clk),
    .D(net912),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7653_ (.CLK(clknet_leaf_89_clk),
    .D(net908),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7654_ (.CLK(clknet_leaf_84_clk),
    .D(net671),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7655_ (.CLK(clknet_leaf_75_clk),
    .D(net669),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7656_ (.CLK(clknet_leaf_75_clk),
    .D(net673),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7657_ (.CLK(clknet_leaf_74_clk),
    .D(net1099),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7658_ (.CLK(clknet_leaf_79_clk),
    .D(net934),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7659_ (.CLK(clknet_leaf_78_clk),
    .D(net1311),
    .Q(\U_DATAPATH.U_ID_EX.o_pc_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7660_ (.CLK(clknet_leaf_48_clk),
    .D(_0636_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7661_ (.CLK(clknet_leaf_48_clk),
    .D(_0637_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7662_ (.CLK(clknet_leaf_55_clk),
    .D(_0638_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7663_ (.CLK(clknet_leaf_55_clk),
    .D(_0639_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7664_ (.CLK(clknet_leaf_53_clk),
    .D(_0640_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7665_ (.CLK(clknet_leaf_53_clk),
    .D(_0641_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7666_ (.CLK(clknet_leaf_51_clk),
    .D(_0642_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7667_ (.CLK(clknet_leaf_50_clk),
    .D(_0643_),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7668_ (.CLK(clknet_leaf_48_clk),
    .D(_0644_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7669_ (.CLK(clknet_leaf_48_clk),
    .D(_0645_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7670_ (.CLK(clknet_leaf_43_clk),
    .D(_0646_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7671_ (.CLK(clknet_leaf_43_clk),
    .D(_0647_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7672_ (.CLK(clknet_leaf_96_clk),
    .D(_0648_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7673_ (.CLK(clknet_leaf_17_clk),
    .D(_0649_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7674_ (.CLK(clknet_leaf_26_clk),
    .D(_0650_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7675_ (.CLK(clknet_leaf_101_clk),
    .D(_0651_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7676_ (.CLK(clknet_leaf_46_clk),
    .D(_0652_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7677_ (.CLK(clknet_leaf_42_clk),
    .D(_0653_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7678_ (.CLK(clknet_leaf_40_clk),
    .D(_0654_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7679_ (.CLK(clknet_leaf_8_clk),
    .D(_0655_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7680_ (.CLK(clknet_leaf_42_clk),
    .D(_0656_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7681_ (.CLK(clknet_leaf_43_clk),
    .D(_0657_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7682_ (.CLK(clknet_leaf_15_clk),
    .D(_0658_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7683_ (.CLK(clknet_leaf_2_clk),
    .D(_0659_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7684_ (.CLK(clknet_leaf_12_clk),
    .D(_0660_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7685_ (.CLK(clknet_leaf_49_clk),
    .D(_0661_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7686_ (.CLK(clknet_leaf_106_clk),
    .D(_0662_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7687_ (.CLK(clknet_leaf_8_clk),
    .D(_0663_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7688_ (.CLK(clknet_leaf_104_clk),
    .D(_0664_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7689_ (.CLK(clknet_leaf_19_clk),
    .D(_0665_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7690_ (.CLK(clknet_leaf_102_clk),
    .D(_0666_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7691_ (.CLK(clknet_leaf_96_clk),
    .D(_0667_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7692_ (.CLK(clknet_leaf_96_clk),
    .D(_0668_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7693_ (.CLK(clknet_leaf_12_clk),
    .D(_0669_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7694_ (.CLK(clknet_leaf_106_clk),
    .D(_0670_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7695_ (.CLK(clknet_leaf_96_clk),
    .D(_0671_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7696_ (.CLK(clknet_leaf_13_clk),
    .D(_0672_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7697_ (.CLK(clknet_leaf_100_clk),
    .D(_0673_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7698_ (.CLK(clknet_leaf_11_clk),
    .D(_0674_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7699_ (.CLK(clknet_leaf_13_clk),
    .D(_0675_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs2_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7700_ (.CLK(clknet_leaf_50_clk),
    .D(_0676_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7701_ (.CLK(clknet_leaf_49_clk),
    .D(_0677_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7702_ (.CLK(clknet_leaf_43_clk),
    .D(_0678_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7703_ (.CLK(clknet_leaf_43_clk),
    .D(_0679_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7704_ (.CLK(clknet_leaf_96_clk),
    .D(_0680_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7705_ (.CLK(clknet_leaf_17_clk),
    .D(_0681_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7706_ (.CLK(clknet_leaf_34_clk),
    .D(_0682_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7707_ (.CLK(clknet_leaf_101_clk),
    .D(_0683_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7708_ (.CLK(clknet_leaf_49_clk),
    .D(_0684_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7709_ (.CLK(clknet_leaf_34_clk),
    .D(_0685_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7710_ (.CLK(clknet_leaf_40_clk),
    .D(_0686_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7711_ (.CLK(clknet_leaf_9_clk),
    .D(_0687_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7712_ (.CLK(clknet_leaf_34_clk),
    .D(_0688_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7713_ (.CLK(clknet_leaf_43_clk),
    .D(_0689_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7714_ (.CLK(clknet_leaf_16_clk),
    .D(_0690_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7715_ (.CLK(clknet_leaf_10_clk),
    .D(_0691_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7716_ (.CLK(clknet_leaf_8_clk),
    .D(_0692_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7717_ (.CLK(clknet_leaf_17_clk),
    .D(_0693_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7718_ (.CLK(clknet_leaf_112_clk),
    .D(_0694_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7719_ (.CLK(clknet_leaf_8_clk),
    .D(_0695_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7720_ (.CLK(clknet_leaf_2_clk),
    .D(_0696_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7721_ (.CLK(clknet_leaf_19_clk),
    .D(_0697_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7722_ (.CLK(clknet_leaf_103_clk),
    .D(_0698_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7723_ (.CLK(clknet_leaf_106_clk),
    .D(_0699_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7724_ (.CLK(clknet_leaf_96_clk),
    .D(_0700_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7725_ (.CLK(clknet_leaf_12_clk),
    .D(_0701_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7726_ (.CLK(clknet_leaf_106_clk),
    .D(_0702_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7727_ (.CLK(clknet_leaf_96_clk),
    .D(_0703_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7728_ (.CLK(clknet_leaf_13_clk),
    .D(_0704_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7729_ (.CLK(clknet_leaf_100_clk),
    .D(_0705_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7730_ (.CLK(clknet_leaf_11_clk),
    .D(_0706_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7731_ (.CLK(clknet_leaf_14_clk),
    .D(_0707_),
    .Q(\U_DATAPATH.U_ID_EX.o_rs1_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7732_ (.CLK(clknet_leaf_55_clk),
    .D(_0708_),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7733_ (.CLK(clknet_leaf_53_clk),
    .D(net1992),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7734_ (.CLK(clknet_leaf_53_clk),
    .D(_0710_),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7735_ (.CLK(clknet_leaf_54_clk),
    .D(_0711_),
    .Q(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7736_ (.CLK(clknet_leaf_71_clk),
    .D(_0712_),
    .Q(\U_CONTROL_UNIT.i_branch_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7737_ (.CLK(clknet_leaf_73_clk),
    .D(_0713_),
    .Q(\U_CONTROL_UNIT.i_jump_EX ));
 sky130_fd_sc_hd__dfxtp_1 _7738_ (.CLK(clknet_leaf_47_clk),
    .D(net954),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7739_ (.CLK(clknet_leaf_47_clk),
    .D(net928),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7740_ (.CLK(clknet_leaf_64_clk),
    .D(_0716_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7741_ (.CLK(clknet_leaf_67_clk),
    .D(_0717_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7742_ (.CLK(clknet_leaf_77_clk),
    .D(_0718_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7743_ (.CLK(clknet_leaf_68_clk),
    .D(_0719_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7744_ (.CLK(clknet_leaf_67_clk),
    .D(_0720_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7745_ (.CLK(clknet_leaf_77_clk),
    .D(_0721_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7746_ (.CLK(clknet_leaf_65_clk),
    .D(_0722_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7747_ (.CLK(clknet_leaf_63_clk),
    .D(_0723_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7748_ (.CLK(clknet_leaf_63_clk),
    .D(_0724_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7749_ (.CLK(clknet_leaf_55_clk),
    .D(_0725_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7750_ (.CLK(clknet_leaf_57_clk),
    .D(_0726_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7751_ (.CLK(clknet_leaf_61_clk),
    .D(_0727_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7752_ (.CLK(clknet_leaf_61_clk),
    .D(_0728_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7753_ (.CLK(clknet_leaf_93_clk),
    .D(_0729_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7754_ (.CLK(clknet_leaf_95_clk),
    .D(_0730_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7755_ (.CLK(clknet_leaf_91_clk),
    .D(_0731_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7756_ (.CLK(clknet_leaf_82_clk),
    .D(_0732_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7757_ (.CLK(clknet_leaf_97_clk),
    .D(_0733_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7758_ (.CLK(clknet_leaf_88_clk),
    .D(_0734_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7759_ (.CLK(clknet_leaf_98_clk),
    .D(_0735_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7760_ (.CLK(clknet_leaf_90_clk),
    .D(_0736_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7761_ (.CLK(clknet_leaf_91_clk),
    .D(_0737_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7762_ (.CLK(clknet_leaf_89_clk),
    .D(_0738_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7763_ (.CLK(clknet_leaf_82_clk),
    .D(_0739_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7764_ (.CLK(clknet_leaf_83_clk),
    .D(_0740_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7765_ (.CLK(clknet_leaf_79_clk),
    .D(_0741_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7766_ (.CLK(clknet_leaf_75_clk),
    .D(_0742_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7767_ (.CLK(clknet_leaf_81_clk),
    .D(_0743_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7768_ (.CLK(clknet_leaf_79_clk),
    .D(_0744_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7769_ (.CLK(clknet_leaf_76_clk),
    .D(_0745_),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_target_M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7770_ (.CLK(clknet_leaf_38_clk),
    .D(net918),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7771_ (.CLK(clknet_leaf_38_clk),
    .D(net846),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7772_ (.CLK(clknet_leaf_38_clk),
    .D(net866),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7773_ (.CLK(clknet_leaf_35_clk),
    .D(net1605),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7774_ (.CLK(clknet_leaf_107_clk),
    .D(net1333),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7775_ (.CLK(clknet_leaf_24_clk),
    .D(net1109),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7776_ (.CLK(clknet_leaf_29_clk),
    .D(net998),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7777_ (.CLK(clknet_leaf_103_clk),
    .D(net1535),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7778_ (.CLK(clknet_leaf_40_clk),
    .D(net1257),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7779_ (.CLK(clknet_leaf_28_clk),
    .D(net1119),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7780_ (.CLK(clknet_leaf_33_clk),
    .D(net1391),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7781_ (.CLK(clknet_leaf_4_clk),
    .D(net1371),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7782_ (.CLK(clknet_leaf_32_clk),
    .D(net1217),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7783_ (.CLK(clknet_leaf_17_clk),
    .D(net1759),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7784_ (.CLK(clknet_leaf_21_clk),
    .D(net1261),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7785_ (.CLK(clknet_leaf_4_clk),
    .D(net1063),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7786_ (.CLK(clknet_leaf_22_clk),
    .D(net1385),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7787_ (.CLK(clknet_leaf_26_clk),
    .D(net1491),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7788_ (.CLK(clknet_leaf_113_clk),
    .D(net1101),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7789_ (.CLK(clknet_leaf_5_clk),
    .D(net1345),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7790_ (.CLK(clknet_leaf_116_clk),
    .D(net1071),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7791_ (.CLK(clknet_leaf_23_clk),
    .D(net1289),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7792_ (.CLK(clknet_leaf_104_clk),
    .D(net1711),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7793_ (.CLK(clknet_leaf_113_clk),
    .D(net1145),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7794_ (.CLK(clknet_leaf_108_clk),
    .D(net1679),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7795_ (.CLK(clknet_leaf_7_clk),
    .D(net1485),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7796_ (.CLK(clknet_leaf_110_clk),
    .D(net1113),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7797_ (.CLK(clknet_leaf_109_clk),
    .D(net1367),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7798_ (.CLK(clknet_leaf_8_clk),
    .D(net1437),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7799_ (.CLK(clknet_leaf_107_clk),
    .D(net1681),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7800_ (.CLK(clknet_leaf_2_clk),
    .D(net1553),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7801_ (.CLK(clknet_leaf_15_clk),
    .D(net1295),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7802_ (.CLK(clknet_leaf_39_clk),
    .D(net830),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7803_ (.CLK(clknet_leaf_38_clk),
    .D(net1049),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7804_ (.CLK(clknet_leaf_41_clk),
    .D(net1301),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7805_ (.CLK(clknet_leaf_39_clk),
    .D(net882),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7806_ (.CLK(clknet_leaf_107_clk),
    .D(net1195),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7807_ (.CLK(clknet_leaf_25_clk),
    .D(net1431),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7808_ (.CLK(clknet_leaf_29_clk),
    .D(net1265),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7809_ (.CLK(clknet_leaf_103_clk),
    .D(net1609),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7810_ (.CLK(clknet_leaf_40_clk),
    .D(net1097),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7811_ (.CLK(clknet_leaf_25_clk),
    .D(net1641),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7812_ (.CLK(clknet_leaf_33_clk),
    .D(net1139),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7813_ (.CLK(clknet_leaf_3_clk),
    .D(net1517),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7814_ (.CLK(clknet_leaf_33_clk),
    .D(net1037),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7815_ (.CLK(clknet_leaf_42_clk),
    .D(net1441),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7816_ (.CLK(clknet_leaf_18_clk),
    .D(net1171),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7817_ (.CLK(clknet_leaf_1_clk),
    .D(net1425),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7818_ (.CLK(clknet_leaf_7_clk),
    .D(net1435),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7819_ (.CLK(clknet_leaf_26_clk),
    .D(net1567),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7820_ (.CLK(clknet_leaf_113_clk),
    .D(net1006),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7821_ (.CLK(clknet_leaf_7_clk),
    .D(net1495),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7822_ (.CLK(clknet_leaf_1_clk),
    .D(net1043),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7823_ (.CLK(clknet_leaf_20_clk),
    .D(net1103),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7824_ (.CLK(clknet_leaf_103_clk),
    .D(net1369),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7825_ (.CLK(clknet_leaf_112_clk),
    .D(net1267),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7826_ (.CLK(clknet_leaf_107_clk),
    .D(net1477),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7827_ (.CLK(clknet_leaf_15_clk),
    .D(net1002),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7828_ (.CLK(clknet_leaf_111_clk),
    .D(net960),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7829_ (.CLK(clknet_leaf_105_clk),
    .D(net1493),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7830_ (.CLK(clknet_leaf_11_clk),
    .D(net1219),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7831_ (.CLK(clknet_leaf_106_clk),
    .D(net1211),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7832_ (.CLK(clknet_leaf_10_clk),
    .D(net1315),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7833_ (.CLK(clknet_leaf_16_clk),
    .D(net1277),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7834_ (.CLK(clknet_leaf_55_clk),
    .D(_0810_),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7835_ (.CLK(clknet_leaf_53_clk),
    .D(_0811_),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7836_ (.CLK(clknet_leaf_53_clk),
    .D(_0812_),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7837_ (.CLK(clknet_leaf_55_clk),
    .D(net862),
    .Q(\U_DATAPATH.U_EX_MEM.o_rd_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7838_ (.CLK(clknet_leaf_64_clk),
    .D(net708),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7839_ (.CLK(clknet_leaf_68_clk),
    .D(net720),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7840_ (.CLK(clknet_leaf_79_clk),
    .D(net641),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7841_ (.CLK(clknet_leaf_78_clk),
    .D(net724),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7842_ (.CLK(clknet_leaf_66_clk),
    .D(net722),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7843_ (.CLK(clknet_leaf_69_clk),
    .D(net816),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7844_ (.CLK(clknet_leaf_65_clk),
    .D(net750),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7845_ (.CLK(clknet_leaf_65_clk),
    .D(net754),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7846_ (.CLK(clknet_leaf_62_clk),
    .D(net691),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7847_ (.CLK(clknet_leaf_54_clk),
    .D(net736),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7848_ (.CLK(clknet_leaf_57_clk),
    .D(net732),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7849_ (.CLK(clknet_leaf_60_clk),
    .D(net758),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7850_ (.CLK(clknet_leaf_61_clk),
    .D(net655),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7851_ (.CLK(clknet_leaf_93_clk),
    .D(net683),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7852_ (.CLK(clknet_leaf_93_clk),
    .D(net778),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7853_ (.CLK(clknet_leaf_91_clk),
    .D(net710),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7854_ (.CLK(clknet_leaf_82_clk),
    .D(net808),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7855_ (.CLK(clknet_leaf_98_clk),
    .D(net812),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7856_ (.CLK(clknet_leaf_88_clk),
    .D(net712),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7857_ (.CLK(clknet_leaf_98_clk),
    .D(net623),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7858_ (.CLK(clknet_leaf_88_clk),
    .D(net633),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7859_ (.CLK(clknet_leaf_92_clk),
    .D(net806),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7860_ (.CLK(clknet_leaf_87_clk),
    .D(net728),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7861_ (.CLK(clknet_leaf_81_clk),
    .D(net760),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7862_ (.CLK(clknet_leaf_84_clk),
    .D(net685),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7863_ (.CLK(clknet_leaf_79_clk),
    .D(net756),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7864_ (.CLK(clknet_leaf_77_clk),
    .D(net657),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7865_ (.CLK(clknet_leaf_81_clk),
    .D(net748),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7866_ (.CLK(clknet_leaf_79_clk),
    .D(net782),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7867_ (.CLK(clknet_leaf_76_clk),
    .D(net792),
    .Q(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7868_ (.CLK(clknet_leaf_48_clk),
    .D(net2343),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7869_ (.CLK(clknet_leaf_49_clk),
    .D(_0845_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7870_ (.CLK(clknet_leaf_44_clk),
    .D(_0846_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7871_ (.CLK(clknet_4_9_0_clk),
    .D(_0847_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7872_ (.CLK(clknet_leaf_98_clk),
    .D(_0848_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7873_ (.CLK(clknet_leaf_16_clk),
    .D(_0849_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7874_ (.CLK(clknet_leaf_42_clk),
    .D(net2359),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7875_ (.CLK(clknet_leaf_73_clk),
    .D(_0851_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7876_ (.CLK(clknet_leaf_46_clk),
    .D(net2346),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7877_ (.CLK(clknet_leaf_48_clk),
    .D(_0853_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7878_ (.CLK(clknet_leaf_49_clk),
    .D(net2339),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7879_ (.CLK(clknet_leaf_12_clk),
    .D(_0855_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7880_ (.CLK(clknet_leaf_40_clk),
    .D(net2371),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7881_ (.CLK(clknet_leaf_44_clk),
    .D(net2382),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7882_ (.CLK(clknet_leaf_16_clk),
    .D(net2375),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7883_ (.CLK(clknet_leaf_13_clk),
    .D(_0859_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7884_ (.CLK(clknet_leaf_12_clk),
    .D(net2350),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7885_ (.CLK(clknet_leaf_44_clk),
    .D(_0861_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7886_ (.CLK(clknet_leaf_102_clk),
    .D(_0862_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7887_ (.CLK(clknet_leaf_13_clk),
    .D(net2368),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7888_ (.CLK(clknet_leaf_100_clk),
    .D(_0864_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7889_ (.CLK(clknet_leaf_12_clk),
    .D(net2378),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7890_ (.CLK(clknet_leaf_99_clk),
    .D(_0866_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7891_ (.CLK(clknet_leaf_100_clk),
    .D(net2392),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7892_ (.CLK(clknet_leaf_98_clk),
    .D(_0868_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7893_ (.CLK(clknet_leaf_13_clk),
    .D(_0869_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7894_ (.CLK(clknet_leaf_98_clk),
    .D(_0870_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7895_ (.CLK(clknet_leaf_98_clk),
    .D(_0871_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7896_ (.CLK(clknet_leaf_76_clk),
    .D(_0872_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7897_ (.CLK(clknet_leaf_98_clk),
    .D(_0873_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7898_ (.CLK(clknet_leaf_13_clk),
    .D(_0874_),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7899_ (.CLK(clknet_leaf_73_clk),
    .D(net2355),
    .Q(\U_DATAPATH.U_EX_MEM.o_alu_result_M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7900_ (.CLK(clknet_leaf_56_clk),
    .D(net1343),
    .Q(\U_DATAPATH.U_EX_MEM.o_result_src_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7901_ (.CLK(clknet_leaf_56_clk),
    .D(net1717),
    .Q(\U_DATAPATH.U_EX_MEM.o_result_src_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7902_ (.CLK(clknet_leaf_56_clk),
    .D(net796),
    .Q(\U_DATAPATH.U_EX_MEM.o_reg_write_M ));
 sky130_fd_sc_hd__dfxtp_1 _7903_ (.CLK(clknet_leaf_86_clk),
    .D(_0879_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7904_ (.CLK(clknet_leaf_4_clk),
    .D(net2308),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7905_ (.CLK(clknet_leaf_94_clk),
    .D(_0881_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7906_ (.CLK(clknet_leaf_22_clk),
    .D(_0882_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7907_ (.CLK(clknet_leaf_54_clk),
    .D(_0883_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7908_ (.CLK(clknet_leaf_30_clk),
    .D(_0884_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7909_ (.CLK(clknet_leaf_32_clk),
    .D(_0885_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7910_ (.CLK(clknet_leaf_92_clk),
    .D(_0886_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7911_ (.CLK(clknet_leaf_23_clk),
    .D(_0887_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7912_ (.CLK(clknet_leaf_29_clk),
    .D(_0888_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7913_ (.CLK(clknet_leaf_59_clk),
    .D(_0889_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7914_ (.CLK(clknet_leaf_24_clk),
    .D(_0890_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7915_ (.CLK(clknet_leaf_28_clk),
    .D(_0891_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7916_ (.CLK(clknet_leaf_0_clk),
    .D(_0892_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7917_ (.CLK(clknet_leaf_115_clk),
    .D(_0893_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7918_ (.CLK(clknet_leaf_116_clk),
    .D(_0894_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7919_ (.CLK(clknet_leaf_5_clk),
    .D(_0895_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7920_ (.CLK(clknet_leaf_52_clk),
    .D(net2126),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7921_ (.CLK(clknet_leaf_52_clk),
    .D(_0897_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7922_ (.CLK(clknet_leaf_6_clk),
    .D(_0898_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7923_ (.CLK(clknet_leaf_115_clk),
    .D(_0899_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7924_ (.CLK(clknet_leaf_0_clk),
    .D(_0900_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7925_ (.CLK(clknet_leaf_52_clk),
    .D(_0901_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7926_ (.CLK(clknet_leaf_94_clk),
    .D(_0902_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7927_ (.CLK(clknet_leaf_57_clk),
    .D(_0903_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7928_ (.CLK(clknet_leaf_85_clk),
    .D(_0904_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7929_ (.CLK(clknet_leaf_115_clk),
    .D(_0905_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7930_ (.CLK(clknet_leaf_115_clk),
    .D(_0906_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7931_ (.CLK(clknet_leaf_114_clk),
    .D(_0907_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7932_ (.CLK(clknet_leaf_109_clk),
    .D(_0908_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7933_ (.CLK(clknet_leaf_78_clk),
    .D(_0909_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7934_ (.CLK(clknet_leaf_94_clk),
    .D(_0910_),
    .Q(\U_DATAPATH.U_EX_MEM.o_write_data_M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7935_ (.CLK(clknet_leaf_115_clk),
    .D(_0911_),
    .Q(\U_DATAPATH.U_EX_MEM.o_mem_write_M ));
 sky130_fd_sc_hd__dfxtp_1 _7936_ (.CLK(clknet_leaf_50_clk),
    .D(net1489),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_reg_write_WB ));
 sky130_fd_sc_hd__dfxtp_2 _7937_ (.CLK(clknet_leaf_48_clk),
    .D(net2112),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7938_ (.CLK(clknet_leaf_53_clk),
    .D(net2002),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[1] ));
 sky130_fd_sc_hd__dfxtp_4 _7939_ (.CLK(clknet_leaf_53_clk),
    .D(net2095),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[2] ));
 sky130_fd_sc_hd__dfxtp_4 _7940_ (.CLK(clknet_leaf_55_clk),
    .D(net2107),
    .Q(\U_DATAPATH.U_HAZARD_UNIT.i_rdAddr_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7941_ (.CLK(clknet_leaf_64_clk),
    .D(net681),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7942_ (.CLK(clknet_leaf_68_clk),
    .D(net800),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7943_ (.CLK(clknet_leaf_79_clk),
    .D(net790),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7944_ (.CLK(clknet_leaf_78_clk),
    .D(net752),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7945_ (.CLK(clknet_leaf_66_clk),
    .D(net798),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7946_ (.CLK(clknet_leaf_76_clk),
    .D(net607),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7947_ (.CLK(clknet_leaf_65_clk),
    .D(net706),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7948_ (.CLK(clknet_leaf_65_clk),
    .D(net689),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7949_ (.CLK(clknet_leaf_63_clk),
    .D(net619),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7950_ (.CLK(clknet_leaf_55_clk),
    .D(net613),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7951_ (.CLK(clknet_leaf_59_clk),
    .D(net675),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7952_ (.CLK(clknet_leaf_60_clk),
    .D(net786),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7953_ (.CLK(clknet_leaf_60_clk),
    .D(net617),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7954_ (.CLK(clknet_leaf_92_clk),
    .D(net645),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7955_ (.CLK(clknet_leaf_93_clk),
    .D(net776),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7956_ (.CLK(clknet_leaf_88_clk),
    .D(net621),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7957_ (.CLK(clknet_leaf_82_clk),
    .D(net740),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7958_ (.CLK(clknet_leaf_98_clk),
    .D(net772),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7959_ (.CLK(clknet_leaf_88_clk),
    .D(net698),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7960_ (.CLK(clknet_leaf_99_clk),
    .D(net842),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7961_ (.CLK(clknet_leaf_88_clk),
    .D(net742),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7962_ (.CLK(clknet_leaf_91_clk),
    .D(net679),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7963_ (.CLK(clknet_leaf_89_clk),
    .D(net637),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7964_ (.CLK(clknet_leaf_80_clk),
    .D(net635),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7965_ (.CLK(clknet_leaf_80_clk),
    .D(net639),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7966_ (.CLK(clknet_leaf_79_clk),
    .D(net764),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7967_ (.CLK(clknet_leaf_76_clk),
    .D(net667),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7968_ (.CLK(clknet_leaf_80_clk),
    .D(net631),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7969_ (.CLK(clknet_leaf_79_clk),
    .D(net766),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _7970_ (.CLK(clknet_leaf_69_clk),
    .D(net734),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_plus4_WB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7971_ (.CLK(clknet_leaf_47_clk),
    .D(net788),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7972_ (.CLK(clknet_leaf_47_clk),
    .D(net762),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7973_ (.CLK(clknet_leaf_64_clk),
    .D(net718),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7974_ (.CLK(clknet_leaf_68_clk),
    .D(net651),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7975_ (.CLK(clknet_leaf_77_clk),
    .D(net746),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7976_ (.CLK(clknet_leaf_68_clk),
    .D(net677),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7977_ (.CLK(clknet_leaf_66_clk),
    .D(net609),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7978_ (.CLK(clknet_leaf_77_clk),
    .D(net738),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7979_ (.CLK(clknet_leaf_65_clk),
    .D(net726),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7980_ (.CLK(clknet_leaf_64_clk),
    .D(net700),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7981_ (.CLK(clknet_leaf_63_clk),
    .D(net774),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7982_ (.CLK(clknet_leaf_55_clk),
    .D(net770),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7983_ (.CLK(clknet_leaf_62_clk),
    .D(net702),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7984_ (.CLK(clknet_leaf_60_clk),
    .D(net615),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7985_ (.CLK(clknet_leaf_61_clk),
    .D(net730),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7986_ (.CLK(clknet_leaf_92_clk),
    .D(net643),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7987_ (.CLK(clknet_leaf_93_clk),
    .D(net663),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7988_ (.CLK(clknet_leaf_88_clk),
    .D(net629),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7989_ (.CLK(clknet_leaf_82_clk),
    .D(net716),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7990_ (.CLK(clknet_leaf_96_clk),
    .D(net625),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7991_ (.CLK(clknet_leaf_88_clk),
    .D(net714),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7992_ (.CLK(clknet_leaf_98_clk),
    .D(net826),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7993_ (.CLK(clknet_leaf_91_clk),
    .D(net627),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7994_ (.CLK(clknet_leaf_92_clk),
    .D(net659),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7995_ (.CLK(clknet_leaf_88_clk),
    .D(net665),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7996_ (.CLK(clknet_leaf_81_clk),
    .D(net653),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7997_ (.CLK(clknet_leaf_81_clk),
    .D(net647),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7998_ (.CLK(clknet_leaf_79_clk),
    .D(net794),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7999_ (.CLK(clknet_leaf_75_clk),
    .D(net693),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8000_ (.CLK(clknet_leaf_81_clk),
    .D(net780),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8001_ (.CLK(clknet_leaf_79_clk),
    .D(net768),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8002_ (.CLK(clknet_leaf_70_clk),
    .D(net687),
    .Q(\U_DATAPATH.U_MEM_WB.o_pc_target_WB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8003_ (.CLK(clknet_leaf_60_clk),
    .D(_0979_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[0] ));
 sky130_fd_sc_hd__dfxtp_2 _8004_ (.CLK(clknet_leaf_29_clk),
    .D(_0980_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8005_ (.CLK(clknet_leaf_58_clk),
    .D(_0981_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8006_ (.CLK(clknet_leaf_80_clk),
    .D(_0982_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8007_ (.CLK(clknet_leaf_87_clk),
    .D(_0983_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8008_ (.CLK(clknet_leaf_85_clk),
    .D(_0984_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[5] ));
 sky130_fd_sc_hd__dfxtp_2 _8009_ (.CLK(clknet_leaf_22_clk),
    .D(_0985_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[6] ));
 sky130_fd_sc_hd__dfxtp_4 _8010_ (.CLK(clknet_leaf_115_clk),
    .D(_0986_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8011_ (.CLK(clknet_leaf_59_clk),
    .D(_0987_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[8] ));
 sky130_fd_sc_hd__dfxtp_4 _8012_ (.CLK(clknet_leaf_110_clk),
    .D(_0988_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[9] ));
 sky130_fd_sc_hd__dfxtp_2 _8013_ (.CLK(clknet_leaf_28_clk),
    .D(_0989_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[10] ));
 sky130_fd_sc_hd__dfxtp_2 _8014_ (.CLK(clknet_leaf_31_clk),
    .D(_0990_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8015_ (.CLK(clknet_leaf_60_clk),
    .D(_0991_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8016_ (.CLK(clknet_leaf_60_clk),
    .D(_0992_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8017_ (.CLK(clknet_leaf_61_clk),
    .D(_0993_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8018_ (.CLK(clknet_leaf_93_clk),
    .D(_0994_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8019_ (.CLK(clknet_leaf_93_clk),
    .D(_0995_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8020_ (.CLK(clknet_leaf_88_clk),
    .D(_0996_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8021_ (.CLK(clknet_leaf_80_clk),
    .D(_0997_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[18] ));
 sky130_fd_sc_hd__dfxtp_2 _8022_ (.CLK(clknet_leaf_116_clk),
    .D(_0998_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8023_ (.CLK(clknet_leaf_87_clk),
    .D(_0999_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[20] ));
 sky130_fd_sc_hd__dfxtp_2 _8024_ (.CLK(clknet_leaf_52_clk),
    .D(_1000_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8025_ (.CLK(clknet_leaf_92_clk),
    .D(_1001_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8026_ (.CLK(clknet_leaf_92_clk),
    .D(_1002_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8027_ (.CLK(clknet_leaf_92_clk),
    .D(_1003_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8028_ (.CLK(clknet_leaf_58_clk),
    .D(_1004_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[25] ));
 sky130_fd_sc_hd__dfxtp_4 _8029_ (.CLK(clknet_leaf_30_clk),
    .D(_1005_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8030_ (.CLK(clknet_leaf_79_clk),
    .D(_1006_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[27] ));
 sky130_fd_sc_hd__dfxtp_2 _8031_ (.CLK(clknet_leaf_28_clk),
    .D(_1007_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8032_ (.CLK(clknet_leaf_87_clk),
    .D(_1008_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8033_ (.CLK(clknet_leaf_84_clk),
    .D(_1009_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8034_ (.CLK(clknet_leaf_60_clk),
    .D(_1010_),
    .Q(\U_DATAPATH.U_MEM_WB.o_read_data_WB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8035_ (.CLK(net509),
    .D(_1011_),
    .Q(net127));
 sky130_fd_sc_hd__dfxtp_1 _8036_ (.CLK(net510),
    .D(_1012_),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_1 _8037_ (.CLK(net511),
    .D(_1013_),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_1 _8038_ (.CLK(net512),
    .D(_1014_),
    .Q(net152));
 sky130_fd_sc_hd__dfxtp_1 _8039_ (.CLK(net513),
    .D(_1015_),
    .Q(net153));
 sky130_fd_sc_hd__dfxtp_1 _8040_ (.CLK(net514),
    .D(_1016_),
    .Q(net154));
 sky130_fd_sc_hd__dfxtp_1 _8041_ (.CLK(net515),
    .D(_1017_),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_1 _8042_ (.CLK(net516),
    .D(_1018_),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_1 _8043_ (.CLK(net517),
    .D(_1019_),
    .Q(net157));
 sky130_fd_sc_hd__dfxtp_1 _8044_ (.CLK(net518),
    .D(_1020_),
    .Q(net158));
 sky130_fd_sc_hd__dfxtp_1 _8045_ (.CLK(net519),
    .D(_1021_),
    .Q(net128));
 sky130_fd_sc_hd__dfxtp_1 _8046_ (.CLK(net520),
    .D(_1022_),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_1 _8047_ (.CLK(net521),
    .D(_1023_),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_1 _8048_ (.CLK(net522),
    .D(_1024_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_1 _8049_ (.CLK(net523),
    .D(_1025_),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_1 _8050_ (.CLK(net524),
    .D(_1026_),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_1 _8051_ (.CLK(net525),
    .D(_1027_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_1 _8052_ (.CLK(net526),
    .D(_1028_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_1 _8053_ (.CLK(net527),
    .D(_1029_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_1 _8054_ (.CLK(net528),
    .D(_1030_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_1 _8055_ (.CLK(net529),
    .D(_1031_),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_1 _8056_ (.CLK(net530),
    .D(_1032_),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_1 _8057_ (.CLK(net531),
    .D(_1033_),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_1 _8058_ (.CLK(net532),
    .D(_1034_),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_1 _8059_ (.CLK(net533),
    .D(_1035_),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_1 _8060_ (.CLK(net534),
    .D(_1036_),
    .Q(net144));
 sky130_fd_sc_hd__dfxtp_1 _8061_ (.CLK(net535),
    .D(_1037_),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_1 _8062_ (.CLK(net536),
    .D(_1038_),
    .Q(net146));
 sky130_fd_sc_hd__dfxtp_1 _8063_ (.CLK(net537),
    .D(_1039_),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_1 _8064_ (.CLK(net538),
    .D(_1040_),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_1 _8065_ (.CLK(net539),
    .D(_1041_),
    .Q(net150));
 sky130_fd_sc_hd__dfxtp_1 _8066_ (.CLK(net540),
    .D(_1042_),
    .Q(net151));
 sky130_fd_sc_hd__dfxtp_1 _8067_ (.CLK(clknet_leaf_56_clk),
    .D(net1411),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8068_ (.CLK(clknet_leaf_47_clk),
    .D(_0080_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8069_ (.CLK(clknet_leaf_43_clk),
    .D(net924),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8070_ (.CLK(clknet_leaf_16_clk),
    .D(net611),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8071_ (.CLK(clknet_leaf_82_clk),
    .D(_0095_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8072_ (.CLK(clknet_leaf_17_clk),
    .D(net661),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8073_ (.CLK(clknet_leaf_34_clk),
    .D(net1559),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8074_ (.CLK(clknet_leaf_76_clk),
    .D(_0098_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8075_ (.CLK(clknet_leaf_63_clk),
    .D(_0099_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8076_ (.CLK(clknet_leaf_47_clk),
    .D(_0100_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8077_ (.CLK(clknet_leaf_49_clk),
    .D(_0070_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8078_ (.CLK(clknet_leaf_12_clk),
    .D(_0071_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8079_ (.CLK(clknet_leaf_55_clk),
    .D(_0072_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8080_ (.CLK(clknet_leaf_48_clk),
    .D(_0073_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8081_ (.CLK(clknet_leaf_16_clk),
    .D(_0074_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8082_ (.CLK(clknet_leaf_10_clk),
    .D(_0075_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8083_ (.CLK(clknet_leaf_12_clk),
    .D(_0076_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8084_ (.CLK(clknet_leaf_63_clk),
    .D(_0077_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8085_ (.CLK(clknet_leaf_100_clk),
    .D(net1898),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8086_ (.CLK(clknet_leaf_12_clk),
    .D(_0079_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8087_ (.CLK(clknet_leaf_110_clk),
    .D(_0081_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8088_ (.CLK(clknet_leaf_15_clk),
    .D(_0082_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8089_ (.CLK(clknet_leaf_74_clk),
    .D(_0083_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8090_ (.CLK(clknet_leaf_92_clk),
    .D(_0084_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8091_ (.CLK(clknet_leaf_89_clk),
    .D(_0085_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8092_ (.CLK(clknet_leaf_13_clk),
    .D(_0086_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8093_ (.CLK(clknet_leaf_81_clk),
    .D(_0087_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8094_ (.CLK(clknet_leaf_83_clk),
    .D(_0088_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8095_ (.CLK(clknet_leaf_76_clk),
    .D(_0089_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8096_ (.CLK(clknet_leaf_80_clk),
    .D(_0090_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8097_ (.CLK(clknet_leaf_13_clk),
    .D(_0092_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8098_ (.CLK(clknet_leaf_70_clk),
    .D(_0093_),
    .Q(\U_DATAPATH.U_MEM_WB.o_alu_result_WB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8099_ (.CLK(net541),
    .D(_1043_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _8100_ (.CLK(clknet_leaf_72_clk),
    .D(_1044_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_src_EX ));
 sky130_fd_sc_hd__dfxtp_2 _8101_ (.CLK(net542),
    .D(_0069_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_1 _8102_ (.CLK(net543),
    .D(_0080_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_2 _8103_ (.CLK(net544),
    .D(_0091_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_1 _8104_ (.CLK(net545),
    .D(_0094_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_1 _8105_ (.CLK(net546),
    .D(_0095_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_2 _8106_ (.CLK(net547),
    .D(_0096_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_1 _8107_ (.CLK(net548),
    .D(_0097_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_2 _8108_ (.CLK(net549),
    .D(_0098_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_1 _8109_ (.CLK(net550),
    .D(_0099_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_1 _8110_ (.CLK(net551),
    .D(_0100_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_2 _8111_ (.CLK(net552),
    .D(_0070_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_2 _8112_ (.CLK(net553),
    .D(_0071_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_1 _8113_ (.CLK(net554),
    .D(_0072_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _8114_ (.CLK(net555),
    .D(_0073_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_1 _8115_ (.CLK(net556),
    .D(_0074_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_2 _8116_ (.CLK(net557),
    .D(_0075_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_2 _8117_ (.CLK(net558),
    .D(_0076_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_1 _8118_ (.CLK(net559),
    .D(_0077_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_1 _8119_ (.CLK(net560),
    .D(_0078_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _8120_ (.CLK(net561),
    .D(_0079_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _8121_ (.CLK(net562),
    .D(_0081_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_2 _8122_ (.CLK(net563),
    .D(_0082_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_2 _8123_ (.CLK(net564),
    .D(_0083_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_1 _8124_ (.CLK(net565),
    .D(_0084_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _8125_ (.CLK(net566),
    .D(_0085_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_2 _8126_ (.CLK(net567),
    .D(_0086_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _8127_ (.CLK(net568),
    .D(_0087_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _8128_ (.CLK(net569),
    .D(_0088_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_2 _8129_ (.CLK(net570),
    .D(_0089_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_1 _8130_ (.CLK(net571),
    .D(_0090_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_2 _8131_ (.CLK(net572),
    .D(_0092_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_2 _8132_ (.CLK(net573),
    .D(_0093_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _8133_ (.CLK(clknet_leaf_40_clk),
    .D(net1253),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8134_ (.CLK(clknet_leaf_40_clk),
    .D(net1329),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8135_ (.CLK(clknet_leaf_41_clk),
    .D(net910),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8136_ (.CLK(clknet_leaf_41_clk),
    .D(net886),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8137_ (.CLK(clknet_leaf_106_clk),
    .D(net1669),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8138_ (.CLK(clknet_leaf_18_clk),
    .D(net1701),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8139_ (.CLK(clknet_leaf_27_clk),
    .D(net1547),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8140_ (.CLK(clknet_leaf_101_clk),
    .D(net1335),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8141_ (.CLK(clknet_leaf_44_clk),
    .D(net1010),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8142_ (.CLK(clknet_leaf_26_clk),
    .D(net1671),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8143_ (.CLK(clknet_leaf_34_clk),
    .D(net1443),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8144_ (.CLK(clknet_leaf_9_clk),
    .D(net1457),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8145_ (.CLK(clknet_leaf_35_clk),
    .D(net1543),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8146_ (.CLK(clknet_leaf_43_clk),
    .D(net1751),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8147_ (.CLK(clknet_leaf_16_clk),
    .D(net1287),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8148_ (.CLK(clknet_leaf_2_clk),
    .D(net1621),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8149_ (.CLK(clknet_leaf_20_clk),
    .D(net1449),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8150_ (.CLK(clknet_leaf_42_clk),
    .D(net1587),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8151_ (.CLK(clknet_leaf_2_clk),
    .D(net1593),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8152_ (.CLK(clknet_leaf_7_clk),
    .D(net1657),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8153_ (.CLK(clknet_leaf_1_clk),
    .D(net1633),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8154_ (.CLK(clknet_leaf_18_clk),
    .D(net1549),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8155_ (.CLK(clknet_leaf_11_clk),
    .D(net1709),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8156_ (.CLK(clknet_leaf_112_clk),
    .D(net1475),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8157_ (.CLK(clknet_leaf_106_clk),
    .D(net1597),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8158_ (.CLK(clknet_leaf_19_clk),
    .D(net992),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8159_ (.CLK(clknet_leaf_104_clk),
    .D(net1527),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8160_ (.CLK(clknet_leaf_105_clk),
    .D(net1061),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8161_ (.CLK(clknet_leaf_13_clk),
    .D(net1765),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8162_ (.CLK(clknet_leaf_102_clk),
    .D(net1251),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8163_ (.CLK(clknet_leaf_10_clk),
    .D(net1569),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8164_ (.CLK(clknet_leaf_14_clk),
    .D(net1239),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8165_ (.CLK(clknet_leaf_70_clk),
    .D(_1077_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8166_ (.CLK(clknet_leaf_51_clk),
    .D(net1723),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8167_ (.CLK(clknet_leaf_51_clk),
    .D(net1787),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8168_ (.CLK(clknet_leaf_37_clk),
    .D(net2101),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8169_ (.CLK(clknet_leaf_36_clk),
    .D(net1904),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8170_ (.CLK(clknet_leaf_108_clk),
    .D(net1926),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8171_ (.CLK(clknet_leaf_25_clk),
    .D(net1928),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8172_ (.CLK(clknet_leaf_31_clk),
    .D(net1801),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8173_ (.CLK(clknet_leaf_101_clk),
    .D(net1825),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8174_ (.CLK(clknet_leaf_46_clk),
    .D(net1685),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8175_ (.CLK(clknet_leaf_27_clk),
    .D(net1839),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8176_ (.CLK(clknet_leaf_33_clk),
    .D(net1916),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8177_ (.CLK(clknet_leaf_3_clk),
    .D(net1863),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8178_ (.CLK(clknet_leaf_35_clk),
    .D(net1886),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8179_ (.CLK(clknet_leaf_43_clk),
    .D(net1986),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8180_ (.CLK(clknet_leaf_21_clk),
    .D(net1781),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8181_ (.CLK(clknet_leaf_4_clk),
    .D(net1849),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8182_ (.CLK(clknet_leaf_21_clk),
    .D(net1783),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8183_ (.CLK(clknet_leaf_17_clk),
    .D(net1910),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8184_ (.CLK(clknet_leaf_113_clk),
    .D(net1942),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8185_ (.CLK(clknet_leaf_7_clk),
    .D(net1930),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8186_ (.CLK(clknet_leaf_113_clk),
    .D(net1857),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8187_ (.CLK(clknet_leaf_23_clk),
    .D(net1888),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8188_ (.CLK(clknet_leaf_104_clk),
    .D(net1912),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8189_ (.CLK(clknet_leaf_110_clk),
    .D(net1940),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8190_ (.CLK(clknet_leaf_94_clk),
    .D(net1795),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8191_ (.CLK(clknet_leaf_8_clk),
    .D(net1896),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8192_ (.CLK(clknet_leaf_109_clk),
    .D(net1902),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8193_ (.CLK(clknet_leaf_107_clk),
    .D(net1934),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8194_ (.CLK(clknet_leaf_11_clk),
    .D(net1892),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8195_ (.CLK(clknet_leaf_96_clk),
    .D(net1869),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8196_ (.CLK(clknet_leaf_104_clk),
    .D(net1924),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8197_ (.CLK(clknet_leaf_15_clk),
    .D(net1944),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8198_ (.CLK(clknet_leaf_38_clk),
    .D(net880),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8199_ (.CLK(clknet_leaf_38_clk),
    .D(net1075),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8200_ (.CLK(clknet_leaf_38_clk),
    .D(net858),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8201_ (.CLK(clknet_leaf_35_clk),
    .D(net1135),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8202_ (.CLK(clknet_leaf_107_clk),
    .D(net1297),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8203_ (.CLK(clknet_leaf_23_clk),
    .D(net1363),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8204_ (.CLK(clknet_leaf_31_clk),
    .D(net1023),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8205_ (.CLK(clknet_leaf_102_clk),
    .D(net1531),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8206_ (.CLK(clknet_leaf_44_clk),
    .D(net972),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8207_ (.CLK(clknet_leaf_24_clk),
    .D(net1179),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8208_ (.CLK(clknet_leaf_31_clk),
    .D(net976),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8209_ (.CLK(clknet_leaf_4_clk),
    .D(net1473),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8210_ (.CLK(clknet_leaf_32_clk),
    .D(net948),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8211_ (.CLK(clknet_leaf_16_clk),
    .D(net1057),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8212_ (.CLK(clknet_leaf_21_clk),
    .D(net1065),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8213_ (.CLK(clknet_leaf_4_clk),
    .D(net1511),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8214_ (.CLK(clknet_leaf_21_clk),
    .D(net1313),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8215_ (.CLK(clknet_leaf_25_clk),
    .D(net1461),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8216_ (.CLK(clknet_leaf_113_clk),
    .D(net1445),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8217_ (.CLK(clknet_leaf_5_clk),
    .D(net1193),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8218_ (.CLK(clknet_leaf_1_clk),
    .D(net1081),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8219_ (.CLK(clknet_leaf_23_clk),
    .D(net1291),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8220_ (.CLK(clknet_leaf_104_clk),
    .D(net1237),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8221_ (.CLK(clknet_leaf_111_clk),
    .D(net1133),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8222_ (.CLK(clknet_leaf_108_clk),
    .D(net1067),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8223_ (.CLK(clknet_leaf_8_clk),
    .D(net1409),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8224_ (.CLK(clknet_leaf_111_clk),
    .D(net1177),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8225_ (.CLK(clknet_leaf_109_clk),
    .D(net1577),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8226_ (.CLK(clknet_leaf_8_clk),
    .D(net1175),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8227_ (.CLK(clknet_leaf_107_clk),
    .D(net1625),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8228_ (.CLK(clknet_leaf_104_clk),
    .D(net1659),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8229_ (.CLK(clknet_leaf_14_clk),
    .D(net1447),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8230_ (.CLK(net574),
    .D(_0032_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8231_ (.CLK(net575),
    .D(_0043_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8232_ (.CLK(net576),
    .D(_0054_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8233_ (.CLK(net577),
    .D(_0057_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8234_ (.CLK(net578),
    .D(_0058_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8235_ (.CLK(net579),
    .D(_0059_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8236_ (.CLK(net580),
    .D(_0060_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8237_ (.CLK(net581),
    .D(_0061_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8238_ (.CLK(net582),
    .D(_0062_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8239_ (.CLK(net583),
    .D(_0063_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8240_ (.CLK(net584),
    .D(_0033_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8241_ (.CLK(net585),
    .D(_0034_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8242_ (.CLK(net586),
    .D(_0035_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8243_ (.CLK(net587),
    .D(_0036_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8244_ (.CLK(net588),
    .D(_0037_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8245_ (.CLK(net589),
    .D(_0038_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8246_ (.CLK(net590),
    .D(_0039_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8247_ (.CLK(net591),
    .D(_0040_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8248_ (.CLK(net592),
    .D(_0041_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8249_ (.CLK(net593),
    .D(_0042_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8250_ (.CLK(net594),
    .D(_0044_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8251_ (.CLK(net595),
    .D(_0045_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8252_ (.CLK(net596),
    .D(_0046_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8253_ (.CLK(net597),
    .D(_0047_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8254_ (.CLK(net598),
    .D(_0048_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8255_ (.CLK(net599),
    .D(_0049_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8256_ (.CLK(net600),
    .D(_0050_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8257_ (.CLK(net601),
    .D(_0051_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8258_ (.CLK(net602),
    .D(_0052_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8259_ (.CLK(net603),
    .D(_0053_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8260_ (.CLK(net604),
    .D(_0055_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8261_ (.CLK(net605),
    .D(_0056_),
    .Q(\U_DATAPATH.U_ID_EX.i_rs1_ID[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8262_ (.CLK(clknet_leaf_38_clk),
    .D(net1373),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8263_ (.CLK(clknet_leaf_37_clk),
    .D(net868),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8264_ (.CLK(clknet_leaf_37_clk),
    .D(net832),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8265_ (.CLK(clknet_leaf_35_clk),
    .D(net1321),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8266_ (.CLK(clknet_leaf_108_clk),
    .D(net1627),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8267_ (.CLK(clknet_leaf_24_clk),
    .D(net1041),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8268_ (.CLK(clknet_leaf_31_clk),
    .D(net1379),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8269_ (.CLK(clknet_leaf_103_clk),
    .D(net1197),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8270_ (.CLK(clknet_leaf_44_clk),
    .D(net1187),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8271_ (.CLK(clknet_leaf_24_clk),
    .D(net1157),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8272_ (.CLK(clknet_leaf_31_clk),
    .D(net1033),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8273_ (.CLK(clknet_leaf_4_clk),
    .D(net1469),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8274_ (.CLK(clknet_leaf_32_clk),
    .D(net1045),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8275_ (.CLK(clknet_leaf_17_clk),
    .D(net1607),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8276_ (.CLK(clknet_leaf_21_clk),
    .D(net1207),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8277_ (.CLK(clknet_leaf_0_clk),
    .D(net1309),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8278_ (.CLK(clknet_leaf_22_clk),
    .D(net1189),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8279_ (.CLK(clknet_leaf_25_clk),
    .D(net1703),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8280_ (.CLK(clknet_leaf_114_clk),
    .D(net1231),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8281_ (.CLK(clknet_leaf_5_clk),
    .D(net1697),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8282_ (.CLK(clknet_leaf_116_clk),
    .D(net1575),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8283_ (.CLK(clknet_leaf_23_clk),
    .D(net1707),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8284_ (.CLK(clknet_leaf_104_clk),
    .D(net1399),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8285_ (.CLK(clknet_leaf_113_clk),
    .D(net1143),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8286_ (.CLK(clknet_leaf_108_clk),
    .D(net1403),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8287_ (.CLK(clknet_leaf_8_clk),
    .D(net1617),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8288_ (.CLK(clknet_leaf_110_clk),
    .D(net1161),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8289_ (.CLK(clknet_leaf_109_clk),
    .D(net1579),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8290_ (.CLK(clknet_leaf_8_clk),
    .D(net1377),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8291_ (.CLK(clknet_leaf_107_clk),
    .D(net1259),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8292_ (.CLK(clknet_leaf_2_clk),
    .D(net1361),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8293_ (.CLK(clknet_leaf_15_clk),
    .D(net1241),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8294_ (.CLK(clknet_leaf_53_clk),
    .D(net904),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8295_ (.CLK(clknet_leaf_53_clk),
    .D(net848),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8296_ (.CLK(clknet_leaf_36_clk),
    .D(net1089),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8297_ (.CLK(clknet_leaf_35_clk),
    .D(net1497),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8298_ (.CLK(clknet_leaf_108_clk),
    .D(net1039),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8299_ (.CLK(clknet_leaf_24_clk),
    .D(net1269),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8300_ (.CLK(clknet_leaf_29_clk),
    .D(net1031),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8301_ (.CLK(clknet_leaf_102_clk),
    .D(net1423),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8302_ (.CLK(clknet_leaf_40_clk),
    .D(net1191),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8303_ (.CLK(clknet_leaf_28_clk),
    .D(net1339),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8304_ (.CLK(clknet_leaf_31_clk),
    .D(net1225),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8305_ (.CLK(clknet_leaf_4_clk),
    .D(net1181),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8306_ (.CLK(clknet_leaf_32_clk),
    .D(net1012),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8307_ (.CLK(clknet_leaf_16_clk),
    .D(net1451),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8308_ (.CLK(clknet_leaf_22_clk),
    .D(net1091),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8309_ (.CLK(clknet_leaf_0_clk),
    .D(net1281),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8310_ (.CLK(clknet_leaf_6_clk),
    .D(net1115),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8311_ (.CLK(clknet_leaf_17_clk),
    .D(net1249),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8312_ (.CLK(clknet_leaf_114_clk),
    .D(net1459),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8313_ (.CLK(clknet_leaf_5_clk),
    .D(net1487),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8314_ (.CLK(clknet_leaf_116_clk),
    .D(net984),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8315_ (.CLK(clknet_leaf_22_clk),
    .D(net1051),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8316_ (.CLK(clknet_leaf_103_clk),
    .D(net1263),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8317_ (.CLK(clknet_leaf_114_clk),
    .D(net1205),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8318_ (.CLK(clknet_leaf_108_clk),
    .D(net1545),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8319_ (.CLK(clknet_leaf_8_clk),
    .D(net1083),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8320_ (.CLK(clknet_leaf_109_clk),
    .D(net1539),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8321_ (.CLK(clknet_leaf_109_clk),
    .D(net1401),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8322_ (.CLK(clknet_leaf_9_clk),
    .D(net1405),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8323_ (.CLK(clknet_leaf_107_clk),
    .D(net1665),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8324_ (.CLK(clknet_leaf_2_clk),
    .D(net1673),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8325_ (.CLK(clknet_leaf_14_clk),
    .D(net1223),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8326_ (.CLK(clknet_leaf_38_clk),
    .D(net1729),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8327_ (.CLK(clknet_leaf_51_clk),
    .D(net1727),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8328_ (.CLK(clknet_leaf_43_clk),
    .D(net1979),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8329_ (.CLK(clknet_leaf_37_clk),
    .D(net2120),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8330_ (.CLK(clknet_leaf_107_clk),
    .D(net1908),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8331_ (.CLK(clknet_leaf_25_clk),
    .D(net1964),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8332_ (.CLK(clknet_leaf_33_clk),
    .D(net1954),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8333_ (.CLK(clknet_leaf_103_clk),
    .D(net1946),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8334_ (.CLK(clknet_leaf_40_clk),
    .D(net1809),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8335_ (.CLK(clknet_leaf_26_clk),
    .D(net1968),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8336_ (.CLK(clknet_leaf_32_clk),
    .D(net1936),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8337_ (.CLK(clknet_leaf_3_clk),
    .D(net1956),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8338_ (.CLK(clknet_leaf_35_clk),
    .D(net1851),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8339_ (.CLK(clknet_leaf_42_clk),
    .D(net1922),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8340_ (.CLK(clknet_leaf_19_clk),
    .D(net1743),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8341_ (.CLK(clknet_leaf_2_clk),
    .D(net1960),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8342_ (.CLK(clknet_leaf_7_clk),
    .D(net1950),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8343_ (.CLK(clknet_leaf_26_clk),
    .D(net1966),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8344_ (.CLK(clknet_leaf_113_clk),
    .D(net1948),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8345_ (.CLK(clknet_leaf_9_clk),
    .D(net1900),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8346_ (.CLK(clknet_leaf_113_clk),
    .D(net1875),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8347_ (.CLK(clknet_leaf_20_clk),
    .D(net1861),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8348_ (.CLK(clknet_leaf_104_clk),
    .D(net1767),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8349_ (.CLK(clknet_leaf_111_clk),
    .D(net1775),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8350_ (.CLK(clknet_leaf_107_clk),
    .D(net1859),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8351_ (.CLK(clknet_leaf_15_clk),
    .D(net1747),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8352_ (.CLK(clknet_leaf_111_clk),
    .D(net1938),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8353_ (.CLK(clknet_leaf_111_clk),
    .D(net1797),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8354_ (.CLK(clknet_leaf_11_clk),
    .D(net1932),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8355_ (.CLK(clknet_leaf_106_clk),
    .D(net1952),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8356_ (.CLK(clknet_leaf_2_clk),
    .D(net1884),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8357_ (.CLK(clknet_leaf_14_clk),
    .D(net1813),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ));
 sky130_fd_sc_hd__dfstp_1 _8358_ (.CLK(clknet_leaf_71_clk),
    .D(_1238_),
    .SET_B(_0260_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8359_ (.CLK(clknet_leaf_68_clk),
    .D(_1239_),
    .RESET_B(_0261_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8360_ (.CLK(clknet_leaf_78_clk),
    .D(_1240_),
    .RESET_B(_0262_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8361_ (.CLK(clknet_leaf_68_clk),
    .D(_1241_),
    .RESET_B(_0263_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8362_ (.CLK(clknet_leaf_67_clk),
    .D(_1242_),
    .RESET_B(_0264_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8363_ (.CLK(clknet_leaf_69_clk),
    .D(_1243_),
    .RESET_B(_0265_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8364_ (.CLK(clknet_leaf_64_clk),
    .D(_1244_),
    .RESET_B(_0266_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8365_ (.CLK(clknet_leaf_65_clk),
    .D(_1245_),
    .RESET_B(_0267_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8366_ (.CLK(clknet_leaf_62_clk),
    .D(net1995),
    .RESET_B(_0268_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8367_ (.CLK(clknet_leaf_57_clk),
    .D(_1247_),
    .RESET_B(_0269_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8368_ (.CLK(clknet_leaf_57_clk),
    .D(_1248_),
    .RESET_B(_0270_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8369_ (.CLK(clknet_leaf_62_clk),
    .D(_1249_),
    .RESET_B(_0271_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8370_ (.CLK(clknet_leaf_61_clk),
    .D(_1250_),
    .RESET_B(_0272_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8371_ (.CLK(clknet_leaf_95_clk),
    .D(_1251_),
    .RESET_B(_0273_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8372_ (.CLK(clknet_leaf_95_clk),
    .D(_1252_),
    .RESET_B(_0274_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8373_ (.CLK(clknet_leaf_97_clk),
    .D(_1253_),
    .RESET_B(_0275_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8374_ (.CLK(clknet_leaf_90_clk),
    .D(_1254_),
    .RESET_B(_0276_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8375_ (.CLK(clknet_leaf_90_clk),
    .D(_1255_),
    .RESET_B(_0277_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[19] ));
 sky130_fd_sc_hd__dfrtp_1 _8376_ (.CLK(clknet_leaf_90_clk),
    .D(_1256_),
    .RESET_B(_0278_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[20] ));
 sky130_fd_sc_hd__dfrtp_1 _8377_ (.CLK(clknet_leaf_90_clk),
    .D(_1257_),
    .RESET_B(_0279_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8378_ (.CLK(clknet_leaf_90_clk),
    .D(_1258_),
    .RESET_B(_0280_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8379_ (.CLK(clknet_leaf_91_clk),
    .D(net2039),
    .RESET_B(_0281_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8380_ (.CLK(clknet_leaf_83_clk),
    .D(_1260_),
    .RESET_B(_0282_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8381_ (.CLK(clknet_leaf_83_clk),
    .D(_1261_),
    .RESET_B(_0283_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[25] ));
 sky130_fd_sc_hd__dfrtp_1 _8382_ (.CLK(clknet_leaf_83_clk),
    .D(_1262_),
    .RESET_B(_0284_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8383_ (.CLK(clknet_leaf_81_clk),
    .D(_1263_),
    .RESET_B(_0285_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[27] ));
 sky130_fd_sc_hd__dfrtp_1 _8384_ (.CLK(clknet_leaf_77_clk),
    .D(_1264_),
    .RESET_B(_0286_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[28] ));
 sky130_fd_sc_hd__dfrtp_1 _8385_ (.CLK(clknet_leaf_81_clk),
    .D(_1265_),
    .RESET_B(_0287_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[29] ));
 sky130_fd_sc_hd__dfrtp_1 _8386_ (.CLK(clknet_leaf_77_clk),
    .D(_1266_),
    .RESET_B(_0288_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[30] ));
 sky130_fd_sc_hd__dfrtp_1 _8387_ (.CLK(clknet_leaf_77_clk),
    .D(_1267_),
    .RESET_B(_0289_),
    .Q(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8388_ (.CLK(clknet_leaf_50_clk),
    .D(net2135),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8389_ (.CLK(clknet_leaf_51_clk),
    .D(net1761),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8390_ (.CLK(clknet_leaf_36_clk),
    .D(net1695),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8391_ (.CLK(clknet_leaf_36_clk),
    .D(net1918),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8392_ (.CLK(clknet_leaf_94_clk),
    .D(net1882),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8393_ (.CLK(clknet_leaf_24_clk),
    .D(net1741),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8394_ (.CLK(clknet_leaf_29_clk),
    .D(net1771),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8395_ (.CLK(clknet_leaf_100_clk),
    .D(net1753),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8396_ (.CLK(clknet_leaf_49_clk),
    .D(net1855),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8397_ (.CLK(clknet_leaf_28_clk),
    .D(net1789),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8398_ (.CLK(clknet_leaf_32_clk),
    .D(net1827),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8399_ (.CLK(clknet_leaf_5_clk),
    .D(net1769),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8400_ (.CLK(clknet_leaf_36_clk),
    .D(net1805),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8401_ (.CLK(clknet_leaf_16_clk),
    .D(net1779),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8402_ (.CLK(clknet_leaf_21_clk),
    .D(net1721),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8403_ (.CLK(clknet_leaf_0_clk),
    .D(net1845),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8404_ (.CLK(clknet_leaf_6_clk),
    .D(net1749),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8405_ (.CLK(clknet_leaf_17_clk),
    .D(net1977),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8406_ (.CLK(clknet_leaf_114_clk),
    .D(net1831),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8407_ (.CLK(clknet_leaf_5_clk),
    .D(net1763),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8408_ (.CLK(clknet_leaf_114_clk),
    .D(net1799),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8409_ (.CLK(clknet_leaf_22_clk),
    .D(net1865),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8410_ (.CLK(clknet_leaf_102_clk),
    .D(net1815),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8411_ (.CLK(clknet_leaf_110_clk),
    .D(net1733),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8412_ (.CLK(clknet_leaf_94_clk),
    .D(net1843),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8413_ (.CLK(clknet_leaf_20_clk),
    .D(net1739),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8414_ (.CLK(clknet_leaf_109_clk),
    .D(net1871),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8415_ (.CLK(clknet_leaf_109_clk),
    .D(net1803),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8416_ (.CLK(clknet_leaf_9_clk),
    .D(net1823),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8417_ (.CLK(clknet_leaf_95_clk),
    .D(net1715),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8418_ (.CLK(clknet_leaf_2_clk),
    .D(net1837),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8419_ (.CLK(clknet_leaf_13_clk),
    .D(net1841),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8420_ (.CLK(clknet_leaf_51_clk),
    .D(net1705),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8421_ (.CLK(clknet_leaf_51_clk),
    .D(net2124),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8422_ (.CLK(clknet_leaf_36_clk),
    .D(net1735),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8423_ (.CLK(clknet_leaf_36_clk),
    .D(net1819),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8424_ (.CLK(clknet_leaf_109_clk),
    .D(net1811),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8425_ (.CLK(clknet_leaf_24_clk),
    .D(net2169),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8426_ (.CLK(clknet_leaf_29_clk),
    .D(net1745),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8427_ (.CLK(clknet_leaf_102_clk),
    .D(net1719),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8428_ (.CLK(clknet_leaf_40_clk),
    .D(net1737),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8429_ (.CLK(clknet_leaf_28_clk),
    .D(net1757),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8430_ (.CLK(clknet_leaf_31_clk),
    .D(net1877),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8431_ (.CLK(clknet_leaf_4_clk),
    .D(net1791),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8432_ (.CLK(clknet_leaf_32_clk),
    .D(net1829),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8433_ (.CLK(clknet_leaf_16_clk),
    .D(net1873),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8434_ (.CLK(clknet_leaf_22_clk),
    .D(net1906),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8435_ (.CLK(clknet_leaf_0_clk),
    .D(net1835),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8436_ (.CLK(clknet_leaf_6_clk),
    .D(net1853),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8437_ (.CLK(clknet_leaf_17_clk),
    .D(net2157),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8438_ (.CLK(clknet_leaf_114_clk),
    .D(net1847),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8439_ (.CLK(clknet_leaf_5_clk),
    .D(net1975),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8440_ (.CLK(clknet_leaf_116_clk),
    .D(net1731),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8441_ (.CLK(clknet_leaf_22_clk),
    .D(net1725),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8442_ (.CLK(clknet_leaf_104_clk),
    .D(net1833),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8443_ (.CLK(clknet_leaf_114_clk),
    .D(net1914),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8444_ (.CLK(clknet_leaf_94_clk),
    .D(net1807),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8445_ (.CLK(clknet_leaf_7_clk),
    .D(net1890),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8446_ (.CLK(clknet_leaf_110_clk),
    .D(net1755),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8447_ (.CLK(clknet_leaf_109_clk),
    .D(net1920),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8448_ (.CLK(clknet_leaf_9_clk),
    .D(net1962),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8449_ (.CLK(clknet_leaf_95_clk),
    .D(net1777),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8450_ (.CLK(clknet_leaf_2_clk),
    .D(net1867),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8451_ (.CLK(clknet_leaf_15_clk),
    .D(net1817),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8452_ (.CLK(clknet_leaf_56_clk),
    .D(_1332_),
    .Q(\U_DATAPATH.U_EX_MEM.i_result_src_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8453_ (.CLK(clknet_leaf_70_clk),
    .D(_1333_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8454_ (.CLK(clknet_leaf_73_clk),
    .D(_1334_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8455_ (.CLK(clknet_leaf_70_clk),
    .D(_1335_),
    .Q(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8456_ (.CLK(clknet_leaf_53_clk),
    .D(net1615),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8457_ (.CLK(clknet_leaf_52_clk),
    .D(net1499),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8458_ (.CLK(clknet_leaf_37_clk),
    .D(net1185),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8459_ (.CLK(clknet_leaf_36_clk),
    .D(net1687),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8460_ (.CLK(clknet_leaf_108_clk),
    .D(net1327),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8461_ (.CLK(clknet_leaf_25_clk),
    .D(net1653),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8462_ (.CLK(clknet_leaf_31_clk),
    .D(net1303),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8463_ (.CLK(clknet_leaf_100_clk),
    .D(net1293),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8464_ (.CLK(clknet_leaf_49_clk),
    .D(net1337),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8465_ (.CLK(clknet_leaf_28_clk),
    .D(net1677),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8466_ (.CLK(clknet_leaf_32_clk),
    .D(net1325),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8467_ (.CLK(clknet_leaf_3_clk),
    .D(net1611),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8468_ (.CLK(clknet_leaf_36_clk),
    .D(net1557),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8469_ (.CLK(clknet_leaf_16_clk),
    .D(net1483),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8470_ (.CLK(clknet_leaf_22_clk),
    .D(net1349),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8471_ (.CLK(clknet_leaf_0_clk),
    .D(net1599),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8472_ (.CLK(clknet_leaf_6_clk),
    .D(net1433),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8473_ (.CLK(clknet_leaf_17_clk),
    .D(net1649),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8474_ (.CLK(clknet_leaf_114_clk),
    .D(net1519),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8475_ (.CLK(clknet_leaf_5_clk),
    .D(net1613),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8476_ (.CLK(clknet_leaf_114_clk),
    .D(net1637),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8477_ (.CLK(clknet_leaf_22_clk),
    .D(net1629),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8478_ (.CLK(clknet_leaf_103_clk),
    .D(net1515),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8479_ (.CLK(clknet_leaf_110_clk),
    .D(net1347),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8480_ (.CLK(clknet_leaf_94_clk),
    .D(net1693),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8481_ (.CLK(clknet_leaf_19_clk),
    .D(net1541),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8482_ (.CLK(clknet_leaf_109_clk),
    .D(net1453),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8483_ (.CLK(clknet_leaf_109_clk),
    .D(net1619),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8484_ (.CLK(clknet_leaf_10_clk),
    .D(net1675),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8485_ (.CLK(clknet_leaf_95_clk),
    .D(net1501),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8486_ (.CLK(clknet_leaf_112_clk),
    .D(net1509),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8487_ (.CLK(clknet_leaf_14_clk),
    .D(net1589),
    .Q(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8488_ (.CLK(clknet_leaf_76_clk),
    .D(net2091),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8489_ (.CLK(clknet_leaf_76_clk),
    .D(net2050),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8490_ (.CLK(clknet_leaf_74_clk),
    .D(net1973),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8491_ (.CLK(clknet_leaf_75_clk),
    .D(_1371_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8492_ (.CLK(clknet_leaf_75_clk),
    .D(net1880),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8493_ (.CLK(clknet_leaf_74_clk),
    .D(_1373_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8494_ (.CLK(clknet_leaf_75_clk),
    .D(net2085),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8495_ (.CLK(clknet_leaf_74_clk),
    .D(_1375_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8496_ (.CLK(clknet_leaf_74_clk),
    .D(_1376_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8497_ (.CLK(clknet_leaf_74_clk),
    .D(_1377_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8498_ (.CLK(clknet_leaf_74_clk),
    .D(_1378_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8499_ (.CLK(clknet_leaf_74_clk),
    .D(_1379_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8500_ (.CLK(clknet_leaf_76_clk),
    .D(net696),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8501_ (.CLK(clknet_leaf_74_clk),
    .D(_1381_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8502_ (.CLK(clknet_leaf_99_clk),
    .D(_1382_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8503_ (.CLK(clknet_leaf_99_clk),
    .D(_1383_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8504_ (.CLK(clknet_leaf_98_clk),
    .D(_1384_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ));
 sky130_fd_sc_hd__dfxtp_2 _8505_ (.CLK(clknet_leaf_72_clk),
    .D(net2147),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8506_ (.CLK(clknet_leaf_72_clk),
    .D(net1982),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8507_ (.CLK(clknet_leaf_56_clk),
    .D(net2129),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8508_ (.CLK(clknet_leaf_47_clk),
    .D(_1388_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8509_ (.CLK(clknet_leaf_63_clk),
    .D(_1389_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8510_ (.CLK(clknet_leaf_63_clk),
    .D(_1390_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8511_ (.CLK(clknet_leaf_72_clk),
    .D(_1391_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8512_ (.CLK(clknet_leaf_70_clk),
    .D(_1392_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8513_ (.CLK(clknet_leaf_72_clk),
    .D(_1393_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8514_ (.CLK(clknet_leaf_70_clk),
    .D(_1394_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8515_ (.CLK(clknet_leaf_70_clk),
    .D(_1395_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8516_ (.CLK(clknet_leaf_47_clk),
    .D(net2183),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8517_ (.CLK(clknet_leaf_46_clk),
    .D(_1397_),
    .Q(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8518_ (.CLK(clknet_leaf_47_clk),
    .D(_1398_),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_target_EX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8519_ (.CLK(clknet_leaf_47_clk),
    .D(_1399_),
    .Q(\U_DATAPATH.U_EX_MEM.i_pc_target_EX[0] ));
 sky130_fd_sc_hd__ebufn_1 _8527_ (.A(net475),
    .TE_B(_3636_),
    .Z(_0064_));
 sky130_fd_sc_hd__conb_1 _8527__475 (.HI(net475));
 sky130_fd_sc_hd__ebufn_1 _8528_ (.A(net476),
    .TE_B(_3637_),
    .Z(_0065_));
 sky130_fd_sc_hd__conb_1 _8528__476 (.HI(net476));
 sky130_fd_sc_hd__ebufn_1 _8529_ (.A(net470),
    .TE_B(_3638_),
    .Z(_0066_));
 sky130_fd_sc_hd__conb_1 _8529__470 (.LO(net470));
 sky130_fd_sc_hd__ebufn_1 _8530_ (.A(net471),
    .TE_B(_3639_),
    .Z(_0067_));
 sky130_fd_sc_hd__conb_1 _8530__471 (.LO(net471));
 sky130_fd_sc_hd__ebufn_1 _8531_ (.A(net472),
    .TE_B(_3640_),
    .Z(_0068_));
 sky130_fd_sc_hd__conb_1 _8531__472 (.LO(net472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__conb_1 core_473 (.LO(net473));
 sky130_fd_sc_hd__conb_1 core_474 (.LO(net474));
 sky130_fd_sc_hd__buf_4 fanout159 (.A(_2680_),
    .X(net159));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(_2680_),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_8 fanout161 (.A(net163),
    .X(net161));
 sky130_fd_sc_hd__buf_4 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_8 fanout163 (.A(_2562_),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_8 fanout164 (.A(net166),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_8 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_6 fanout166 (.A(_2562_),
    .X(net166));
 sky130_fd_sc_hd__buf_4 fanout167 (.A(net2115),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(net2115),
    .X(net168));
 sky130_fd_sc_hd__buf_4 fanout169 (.A(net173),
    .X(net169));
 sky130_fd_sc_hd__buf_2 fanout170 (.A(net173),
    .X(net170));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(net173),
    .X(net171));
 sky130_fd_sc_hd__buf_4 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(net2115),
    .X(net173));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net2115),
    .X(net174));
 sky130_fd_sc_hd__buf_2 fanout175 (.A(net2115),
    .X(net175));
 sky130_fd_sc_hd__buf_4 fanout176 (.A(net179),
    .X(net176));
 sky130_fd_sc_hd__buf_4 fanout177 (.A(net179),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__buf_6 fanout179 (.A(net2115),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_8 fanout180 (.A(net182),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_8 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(_1722_),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_8 fanout183 (.A(_1721_),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_8 fanout184 (.A(_1721_),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_8 fanout185 (.A(net187),
    .X(net185));
 sky130_fd_sc_hd__buf_4 fanout186 (.A(net187),
    .X(net186));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(_1698_),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_8 fanout188 (.A(_1697_),
    .X(net188));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(_1697_),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_8 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_8 fanout191 (.A(_1681_),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_8 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__buf_6 fanout193 (.A(_1680_),
    .X(net193));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_4 fanout195 (.A(net197),
    .X(net195));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 fanout197 (.A(_1672_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_8 fanout198 (.A(net200),
    .X(net198));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_4 fanout200 (.A(_1671_),
    .X(net200));
 sky130_fd_sc_hd__buf_4 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(_1659_),
    .X(net202));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(_1659_),
    .X(net203));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__buf_4 fanout205 (.A(net207),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_8 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 fanout207 (.A(_1658_),
    .X(net207));
 sky130_fd_sc_hd__buf_4 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_8 fanout209 (.A(_2772_),
    .X(net209));
 sky130_fd_sc_hd__buf_4 fanout210 (.A(_2772_),
    .X(net210));
 sky130_fd_sc_hd__buf_4 fanout211 (.A(_2772_),
    .X(net211));
 sky130_fd_sc_hd__buf_4 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_8 fanout213 (.A(net232),
    .X(net213));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(net219),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_2 fanout215 (.A(net219),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_4 fanout216 (.A(net219),
    .X(net216));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__buf_4 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_4 fanout219 (.A(net232),
    .X(net219));
 sky130_fd_sc_hd__buf_4 fanout220 (.A(net222),
    .X(net220));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 fanout222 (.A(net232),
    .X(net222));
 sky130_fd_sc_hd__buf_4 fanout223 (.A(net232),
    .X(net223));
 sky130_fd_sc_hd__buf_4 fanout224 (.A(net232),
    .X(net224));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(net227),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 fanout226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__buf_4 fanout227 (.A(net232),
    .X(net227));
 sky130_fd_sc_hd__buf_4 fanout228 (.A(net232),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 fanout229 (.A(net232),
    .X(net229));
 sky130_fd_sc_hd__buf_4 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__buf_6 fanout232 (.A(_2122_),
    .X(net232));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net237),
    .X(net233));
 sky130_fd_sc_hd__buf_2 fanout234 (.A(net237),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_8 fanout235 (.A(net237),
    .X(net235));
 sky130_fd_sc_hd__buf_4 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__buf_4 fanout237 (.A(net242),
    .X(net237));
 sky130_fd_sc_hd__buf_4 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 fanout239 (.A(net242),
    .X(net239));
 sky130_fd_sc_hd__buf_4 fanout240 (.A(net241),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_4 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__buf_12 fanout242 (.A(_2121_),
    .X(net242));
 sky130_fd_sc_hd__buf_8 fanout243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_16 fanout244 (.A(_1428_),
    .X(net244));
 sky130_fd_sc_hd__buf_8 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__buf_8 fanout246 (.A(_3482_),
    .X(net246));
 sky130_fd_sc_hd__buf_8 fanout247 (.A(_3478_),
    .X(net247));
 sky130_fd_sc_hd__buf_6 fanout248 (.A(_3478_),
    .X(net248));
 sky130_fd_sc_hd__buf_8 fanout249 (.A(_3474_),
    .X(net249));
 sky130_fd_sc_hd__buf_6 fanout250 (.A(_3474_),
    .X(net250));
 sky130_fd_sc_hd__buf_6 fanout251 (.A(_3429_),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_8 fanout252 (.A(_3429_),
    .X(net252));
 sky130_fd_sc_hd__buf_6 fanout253 (.A(_2724_),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_8 fanout254 (.A(_2724_),
    .X(net254));
 sky130_fd_sc_hd__buf_8 fanout255 (.A(_2720_),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_8 fanout256 (.A(_2720_),
    .X(net256));
 sky130_fd_sc_hd__buf_6 fanout257 (.A(_2677_),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_8 fanout258 (.A(_2677_),
    .X(net258));
 sky130_fd_sc_hd__buf_6 fanout259 (.A(_2673_),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_8 fanout260 (.A(_2673_),
    .X(net260));
 sky130_fd_sc_hd__buf_6 fanout261 (.A(_2668_),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_8 fanout262 (.A(_2668_),
    .X(net262));
 sky130_fd_sc_hd__buf_6 fanout263 (.A(_2664_),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_8 fanout264 (.A(_2664_),
    .X(net264));
 sky130_fd_sc_hd__buf_6 fanout265 (.A(_2658_),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_8 fanout266 (.A(_2658_),
    .X(net266));
 sky130_fd_sc_hd__buf_6 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__buf_8 fanout268 (.A(_1460_),
    .X(net268));
 sky130_fd_sc_hd__buf_6 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__buf_8 fanout270 (.A(_1458_),
    .X(net270));
 sky130_fd_sc_hd__buf_4 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_8 fanout272 (.A(_1436_),
    .X(net272));
 sky130_fd_sc_hd__buf_8 fanout273 (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__buf_12 fanout274 (.A(_1421_),
    .X(net274));
 sky130_fd_sc_hd__buf_8 fanout275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_16 fanout276 (.A(_3553_),
    .X(net276));
 sky130_fd_sc_hd__buf_6 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__buf_8 fanout278 (.A(_3552_),
    .X(net278));
 sky130_fd_sc_hd__buf_8 fanout279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__buf_12 fanout280 (.A(_3519_),
    .X(net280));
 sky130_fd_sc_hd__buf_6 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_8 fanout282 (.A(_3518_),
    .X(net282));
 sky130_fd_sc_hd__buf_6 fanout283 (.A(_3485_),
    .X(net283));
 sky130_fd_sc_hd__buf_6 fanout284 (.A(_3485_),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_8 fanout285 (.A(_3484_),
    .X(net285));
 sky130_fd_sc_hd__buf_4 fanout286 (.A(_3484_),
    .X(net286));
 sky130_fd_sc_hd__buf_8 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__buf_8 fanout288 (.A(_3480_),
    .X(net288));
 sky130_fd_sc_hd__buf_8 fanout289 (.A(_3476_),
    .X(net289));
 sky130_fd_sc_hd__buf_8 fanout290 (.A(_3476_),
    .X(net290));
 sky130_fd_sc_hd__buf_6 fanout291 (.A(_3472_),
    .X(net291));
 sky130_fd_sc_hd__buf_8 fanout292 (.A(_3472_),
    .X(net292));
 sky130_fd_sc_hd__buf_8 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_16 fanout294 (.A(_3439_),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_8 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__buf_8 fanout296 (.A(_3438_),
    .X(net296));
 sky130_fd_sc_hd__buf_6 fanout297 (.A(_3427_),
    .X(net297));
 sky130_fd_sc_hd__buf_6 fanout298 (.A(_3427_),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_8 fanout299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_8 fanout300 (.A(_2769_),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_8 fanout301 (.A(net302),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_8 fanout302 (.A(net2337),
    .X(net302));
 sky130_fd_sc_hd__buf_6 fanout303 (.A(_2722_),
    .X(net303));
 sky130_fd_sc_hd__buf_6 fanout304 (.A(_2722_),
    .X(net304));
 sky130_fd_sc_hd__buf_8 fanout305 (.A(_2718_),
    .X(net305));
 sky130_fd_sc_hd__buf_6 fanout306 (.A(_2718_),
    .X(net306));
 sky130_fd_sc_hd__buf_6 fanout307 (.A(_2675_),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_8 fanout308 (.A(_2675_),
    .X(net308));
 sky130_fd_sc_hd__buf_8 fanout309 (.A(_2671_),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_8 fanout310 (.A(_2671_),
    .X(net310));
 sky130_fd_sc_hd__buf_8 fanout311 (.A(_2666_),
    .X(net311));
 sky130_fd_sc_hd__buf_6 fanout312 (.A(_2666_),
    .X(net312));
 sky130_fd_sc_hd__buf_6 fanout313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__buf_6 fanout314 (.A(_2662_),
    .X(net314));
 sky130_fd_sc_hd__buf_6 fanout315 (.A(_2656_),
    .X(net315));
 sky130_fd_sc_hd__buf_6 fanout316 (.A(_2656_),
    .X(net316));
 sky130_fd_sc_hd__buf_4 fanout317 (.A(_1832_),
    .X(net317));
 sky130_fd_sc_hd__buf_4 fanout318 (.A(_1821_),
    .X(net318));
 sky130_fd_sc_hd__buf_4 fanout319 (.A(_1809_),
    .X(net319));
 sky130_fd_sc_hd__buf_4 fanout320 (.A(_1800_),
    .X(net320));
 sky130_fd_sc_hd__buf_4 fanout321 (.A(_1787_),
    .X(net321));
 sky130_fd_sc_hd__buf_4 fanout322 (.A(_1776_),
    .X(net322));
 sky130_fd_sc_hd__buf_4 fanout323 (.A(_1763_),
    .X(net323));
 sky130_fd_sc_hd__buf_4 fanout324 (.A(_1752_),
    .X(net324));
 sky130_fd_sc_hd__buf_4 fanout325 (.A(_1740_),
    .X(net325));
 sky130_fd_sc_hd__buf_4 fanout326 (.A(_1729_),
    .X(net326));
 sky130_fd_sc_hd__buf_4 fanout327 (.A(_1717_),
    .X(net327));
 sky130_fd_sc_hd__buf_4 fanout328 (.A(_1706_),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_8 fanout329 (.A(_1665_),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_8 fanout330 (.A(_1652_),
    .X(net330));
 sky130_fd_sc_hd__buf_4 fanout331 (.A(_1638_),
    .X(net331));
 sky130_fd_sc_hd__buf_4 fanout332 (.A(_1627_),
    .X(net332));
 sky130_fd_sc_hd__buf_4 fanout333 (.A(_1614_),
    .X(net333));
 sky130_fd_sc_hd__buf_4 fanout334 (.A(_1603_),
    .X(net334));
 sky130_fd_sc_hd__buf_4 fanout335 (.A(_1578_),
    .X(net335));
 sky130_fd_sc_hd__buf_4 fanout336 (.A(_1566_),
    .X(net336));
 sky130_fd_sc_hd__buf_4 fanout337 (.A(_1555_),
    .X(net337));
 sky130_fd_sc_hd__buf_4 fanout338 (.A(_1543_),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_8 fanout339 (.A(_1531_),
    .X(net339));
 sky130_fd_sc_hd__buf_4 fanout340 (.A(_1519_),
    .X(net340));
 sky130_fd_sc_hd__buf_4 fanout341 (.A(_1506_),
    .X(net341));
 sky130_fd_sc_hd__buf_4 fanout342 (.A(_1492_),
    .X(net342));
 sky130_fd_sc_hd__buf_4 fanout343 (.A(_1480_),
    .X(net343));
 sky130_fd_sc_hd__buf_4 fanout344 (.A(_1469_),
    .X(net344));
 sky130_fd_sc_hd__buf_8 fanout345 (.A(net347),
    .X(net345));
 sky130_fd_sc_hd__buf_4 fanout346 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__buf_4 fanout347 (.A(_1448_),
    .X(net347));
 sky130_fd_sc_hd__buf_4 fanout348 (.A(_1435_),
    .X(net348));
 sky130_fd_sc_hd__buf_4 fanout349 (.A(net350),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_8 fanout350 (.A(_2770_),
    .X(net350));
 sky130_fd_sc_hd__buf_4 fanout351 (.A(_2764_),
    .X(net351));
 sky130_fd_sc_hd__buf_4 fanout352 (.A(_2764_),
    .X(net352));
 sky130_fd_sc_hd__buf_8 fanout353 (.A(_2761_),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_8 fanout354 (.A(_2761_),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_8 fanout356 (.A(_1676_),
    .X(net356));
 sky130_fd_sc_hd__buf_4 fanout357 (.A(_1589_),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_8 fanout358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__buf_8 fanout359 (.A(_1433_),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_8 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__buf_8 fanout361 (.A(_1431_),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_16 fanout362 (.A(_1430_),
    .X(net362));
 sky130_fd_sc_hd__buf_6 fanout363 (.A(_1430_),
    .X(net363));
 sky130_fd_sc_hd__buf_8 fanout364 (.A(_1410_),
    .X(net364));
 sky130_fd_sc_hd__buf_4 fanout365 (.A(_1410_),
    .X(net365));
 sky130_fd_sc_hd__buf_8 fanout366 (.A(net2330),
    .X(net366));
 sky130_fd_sc_hd__buf_4 fanout367 (.A(net2330),
    .X(net367));
 sky130_fd_sc_hd__buf_8 fanout368 (.A(net2181),
    .X(net368));
 sky130_fd_sc_hd__buf_8 fanout369 (.A(net2181),
    .X(net369));
 sky130_fd_sc_hd__buf_8 fanout370 (.A(net372),
    .X(net370));
 sky130_fd_sc_hd__buf_4 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__buf_6 fanout372 (.A(net2242),
    .X(net372));
 sky130_fd_sc_hd__buf_8 fanout373 (.A(net375),
    .X(net373));
 sky130_fd_sc_hd__buf_4 fanout374 (.A(net375),
    .X(net374));
 sky130_fd_sc_hd__buf_6 fanout375 (.A(net2242),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_8 fanout376 (.A(net379),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_4 fanout377 (.A(net379),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_8 fanout378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_4 fanout379 (.A(net386),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_8 fanout380 (.A(net386),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_8 fanout381 (.A(net384),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_8 fanout382 (.A(net384),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_4 fanout383 (.A(net384),
    .X(net383));
 sky130_fd_sc_hd__buf_4 fanout384 (.A(net386),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_8 fanout385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_8 fanout386 (.A(net2238),
    .X(net386));
 sky130_fd_sc_hd__buf_8 fanout387 (.A(net390),
    .X(net387));
 sky130_fd_sc_hd__buf_4 fanout388 (.A(net390),
    .X(net388));
 sky130_fd_sc_hd__buf_8 fanout389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__buf_4 fanout390 (.A(net2246),
    .X(net390));
 sky130_fd_sc_hd__buf_8 fanout391 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ),
    .X(net391));
 sky130_fd_sc_hd__buf_8 fanout392 (.A(net396),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_4 fanout393 (.A(net396),
    .X(net393));
 sky130_fd_sc_hd__buf_8 fanout394 (.A(net396),
    .X(net394));
 sky130_fd_sc_hd__buf_4 fanout395 (.A(net396),
    .X(net395));
 sky130_fd_sc_hd__buf_8 fanout396 (.A(net2246),
    .X(net396));
 sky130_fd_sc_hd__buf_8 fanout397 (.A(net399),
    .X(net397));
 sky130_fd_sc_hd__buf_8 fanout398 (.A(net399),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_8 fanout399 (.A(net2264),
    .X(net399));
 sky130_fd_sc_hd__buf_8 fanout400 (.A(net402),
    .X(net400));
 sky130_fd_sc_hd__buf_4 fanout401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__buf_6 fanout402 (.A(net2351),
    .X(net402));
 sky130_fd_sc_hd__buf_8 fanout403 (.A(net404),
    .X(net403));
 sky130_fd_sc_hd__buf_8 fanout404 (.A(net2351),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_8 fanout405 (.A(net408),
    .X(net405));
 sky130_fd_sc_hd__buf_4 fanout406 (.A(net408),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_8 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__buf_4 fanout408 (.A(net409),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_8 fanout409 (.A(net2334),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_8 fanout410 (.A(net411),
    .X(net410));
 sky130_fd_sc_hd__buf_4 fanout411 (.A(net414),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_8 fanout412 (.A(net414),
    .X(net412));
 sky130_fd_sc_hd__buf_4 fanout413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__buf_6 fanout414 (.A(net2334),
    .X(net414));
 sky130_fd_sc_hd__buf_8 fanout415 (.A(net419),
    .X(net415));
 sky130_fd_sc_hd__buf_4 fanout416 (.A(net419),
    .X(net416));
 sky130_fd_sc_hd__buf_8 fanout417 (.A(net419),
    .X(net417));
 sky130_fd_sc_hd__buf_8 fanout418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__buf_8 fanout419 (.A(net2352),
    .X(net419));
 sky130_fd_sc_hd__buf_8 fanout420 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net420));
 sky130_fd_sc_hd__buf_4 fanout421 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net421));
 sky130_fd_sc_hd__buf_8 fanout422 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net422));
 sky130_fd_sc_hd__buf_4 fanout423 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net423));
 sky130_fd_sc_hd__buf_8 fanout424 (.A(net2352),
    .X(net424));
 sky130_fd_sc_hd__buf_4 fanout425 (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_8 fanout426 (.A(\U_DATAPATH.U_MEM_WB.o_result_src_WB[1] ),
    .X(net426));
 sky130_fd_sc_hd__buf_4 fanout427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__buf_4 fanout428 (.A(net431),
    .X(net428));
 sky130_fd_sc_hd__buf_4 fanout429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_4 fanout430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_4 fanout431 (.A(net460),
    .X(net431));
 sky130_fd_sc_hd__buf_4 fanout432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__buf_4 fanout433 (.A(net460),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_8 fanout434 (.A(net460),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_4 fanout435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_4 fanout436 (.A(net437),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_4 fanout437 (.A(net460),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_4 fanout438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__buf_4 fanout439 (.A(net460),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_4 fanout440 (.A(net442),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_4 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_4 fanout442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_4 fanout443 (.A(net460),
    .X(net443));
 sky130_fd_sc_hd__buf_4 fanout444 (.A(net446),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_4 fanout445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__buf_4 fanout446 (.A(net459),
    .X(net446));
 sky130_fd_sc_hd__buf_4 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_4 fanout448 (.A(net459),
    .X(net448));
 sky130_fd_sc_hd__buf_4 fanout449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__buf_4 fanout450 (.A(net459),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_4 fanout451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_4 fanout452 (.A(net459),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_4 fanout453 (.A(net458),
    .X(net453));
 sky130_fd_sc_hd__buf_4 fanout454 (.A(net458),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_4 fanout455 (.A(net457),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_2 fanout456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__buf_2 fanout457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_4 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_8 fanout459 (.A(net460),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_8 fanout460 (.A(_0101_),
    .X(net460));
 sky130_fd_sc_hd__buf_8 fanout461 (.A(net63),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_4 fanout462 (.A(net63),
    .X(net462));
 sky130_fd_sc_hd__buf_8 fanout463 (.A(net465),
    .X(net463));
 sky130_fd_sc_hd__buf_8 fanout464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_8 fanout465 (.A(net63),
    .X(net465));
 sky130_fd_sc_hd__buf_6 fanout466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__buf_6 fanout467 (.A(net63),
    .X(net467));
 sky130_fd_sc_hd__buf_8 fanout468 (.A(net63),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_8 fanout469 (.A(net63),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[7] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0960_),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[8] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(_0749_),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][13] ),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(_1155_),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][7] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(_0785_),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][11] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(_1347_),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][19] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(_1355_),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][0] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_0923_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(_1336_),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][25] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(_1167_),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][27] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(_1363_),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][15] ),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(_1060_),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][29] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(_0441_),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][29] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[2] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(_1139_),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][4] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(_1146_),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][21] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(_1357_),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][12] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(_0552_),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][20] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(_1065_),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][9] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_0814_),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(_0517_),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][20] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(_1356_),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][7] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(_0419_),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][9] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(_0787_),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][17] ),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(_0493_),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][8] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[17] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(_0548_),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][8] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(_0420_),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][17] ),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(_1353_),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][29] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(_0473_),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][5] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(_1341_),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][4] ),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0829_),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(_0480_),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][19] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(_1064_),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][30] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(_1140_),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][4] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(_0544_),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][29] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(_0505_),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][29] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[20] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(_1203_),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][2] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(_0478_),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][4] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(_1049_),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][9] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(_1054_),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][30] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(_1204_),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][28] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0832_),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(_1364_),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][9] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(_1345_),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][24] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(_0770_),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][29] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(_0775_),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][12] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(_0520_),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][8] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[20] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(_1086_),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][3] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(_1339_),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][4] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(_0416_),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][20] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(_0528_),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][24] ),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(_1360_),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][2] ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0967_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(_1270_),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][19] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(_1161_),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][7] ),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(_0483_),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][5] ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(_1050_),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][17] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(_1159_),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][0] ),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[14] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[18] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(_1300_),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][21] ),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(_1163_),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][22] ),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(_1067_),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][22] ),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(_0768_),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][13] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(_0457_),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][29] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0965_),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(_1297_),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\U_DATAPATH.U_EX_MEM.i_result_src_EX[1] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(_0877_),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][7] ),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(_1307_),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][14] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(_1282_),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][0] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(_1078_),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][21] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[2] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(_1321_),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][1] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(_1207_),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][0] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(_1206_),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][20] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(_1320_),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][23] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(_1291_),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][2] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_0949_),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(_1302_),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][8] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(_1308_),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][25] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(_1293_),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][5] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(_1273_),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][14] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(_1220_),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][6] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[3] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(_1306_),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][25] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(_1231_),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][16] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(_1284_),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][13] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(_1058_),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][7] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(_1275_),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][26] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0815_),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(_1326_),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][9] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(_1309_),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][13] ),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(_0759_),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][1] ),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(_1269_),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][19] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(_1287_),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][28] ),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[6] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(_1073_),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][22] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(_1228_),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][11] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(_1279_),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][6] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(_1274_),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][7] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(_0515_),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][23] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0818_),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(_1229_),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][29] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(_1329_),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][13] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(_1281_),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][14] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(_1092_),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][16] ),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(_1094_),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[19] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[5] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(_0339_),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][1] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(_1079_),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][9] ),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(_1277_),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][11] ),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(_1311_),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[13] ),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(_0333_),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][24] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0817_),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(_1102_),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][27] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(_1233_),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][20] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(_1288_),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][6] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(_1084_),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][27] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(_1295_),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][12] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0929_),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[8] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(_1280_),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][24] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(_1324_),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][8] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(_1214_),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][4] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(_1304_),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][31] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(_1237_),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][22] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_0955_),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(_1290_),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][31] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(_1331_),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][3] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(_1303_),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[22] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(_0342_),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][28] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(_1296_),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][7] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[24] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(_1085_),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][10] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(_1278_),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][12] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(_1312_),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][18] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(_1286_),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][22] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(_1322_),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][15] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0836_),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(_1315_),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][30] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(_1298_),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][9] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(_1087_),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][31] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(_1299_),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][24] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(_1292_),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][15] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[14] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(_1283_),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][18] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(_1318_),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][15] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(_1093_),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][12] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(_1218_),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][16] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(_1316_),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][8] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_0961_),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(_1276_),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][20] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(_1098_),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][24] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(_1230_),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][21] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(_1227_),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][11] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(_1089_),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][21] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[12] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(_1289_),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][30] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(_1330_),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][29] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(_1107_),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][26] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(_1294_),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][13] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(_1313_),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][20] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_0824_),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(_1226_),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][10] ),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(_1310_),
    .X(net1877));
 sky130_fd_sc_hd__clkbuf_2 hold1273 (.A(net2419),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(_3611_),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(_1372_),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][4] ),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(_1272_),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][30] ),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(_1236_),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[31] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][12] ),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(_1090_),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][21] ),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(_1099_),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][25] ),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(_1325_),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][28] ),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(_1106_),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[8] ),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(_0328_),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0946_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][25] ),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(_1103_),
    .X(net1896));
 sky130_fd_sc_hd__buf_1 hold1292 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[18] ),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(_0078_),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][19] ),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(_1225_),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][26] ),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(_1104_),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][3] ),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(_1081_),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[10] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[11] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][14] ),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(_1314_),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][4] ),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(_1210_),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][17] ),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(_1095_),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][22] ),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(_1100_),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][23] ),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(_1323_),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_0823_),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][10] ),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(_1088_),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][3] ),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(_1271_),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][27] ),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(_1327_),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][13] ),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(_1219_),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][30] ),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(_1108_),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[7] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][4] ),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(_1082_),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][5] ),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(_1083_),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][19] ),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(_1097_),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][28] ),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(_1234_),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][27] ),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(_1105_),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_0954_),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][10] ),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(_1216_),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][26] ),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(_1232_),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][23] ),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(_1101_),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][18] ),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(_1096_),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][31] ),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(_1109_),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[18] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][7] ),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(_1213_),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][18] ),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(_1224_),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][16] ),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(_1222_),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][29] ),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(_1235_),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][6] ),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(_1212_),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0933_),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][11] ),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(_1217_),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[0] ),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(_1404_),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][15] ),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(_1221_),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][28] ),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(_1328_),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][5] ),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(_1211_),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[22] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][17] ),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(_1223_),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][9] ),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(_1215_),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[21] ),
    .X(net1969));
 sky130_fd_sc_hd__clkbuf_2 hold1365 (.A(net1488),
    .X(net1970));
 sky130_fd_sc_hd__buf_2 hold1366 (.A(net2116),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(_3609_),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(_1370_),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][19] ),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0937_),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(_1319_),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][17] ),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(_1285_),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][2] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(_1208_),
    .X(net1979));
 sky130_fd_sc_hd__clkbuf_4 hold1375 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[1] ),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(_3626_),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(_1386_),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[30] ),
    .X(net1983));
 sky130_fd_sc_hd__buf_1 hold1379 (.A(net2405),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\U_DATAPATH.U_EX_MEM.o_result_src_M[1] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][13] ),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(_1091_),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[18] ),
    .X(net1987));
 sky130_fd_sc_hd__clkbuf_4 hold1383 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[4] ),
    .X(net1988));
 sky130_fd_sc_hd__buf_4 hold1384 (.A(_2699_),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[31] ),
    .X(net1990));
 sky130_fd_sc_hd__clkbuf_2 hold1386 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[1] ),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(_0709_),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[26] ),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[10] ),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_0291_),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(_1246_),
    .X(net1995));
 sky130_fd_sc_hd__buf_1 hold1391 (.A(net2409),
    .X(net1996));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1392 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[16] ),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[9] ),
    .X(net1998));
 sky130_fd_sc_hd__buf_1 hold1394 (.A(net2111),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[24] ),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[7] ),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(_0914_),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[12] ),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(_1978_),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0925_),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[4] ),
    .X(net745));
 sky130_fd_sc_hd__buf_1 hold1400 (.A(_1979_),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(_2153_),
    .X(net2006));
 sky130_fd_sc_hd__clkbuf_2 hold1402 (.A(net2010),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[29] ),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(_2099_),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[17] ),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[28] ),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[18] ),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(_2016_),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(_2017_),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_0951_),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(_2019_),
    .X(net2015));
 sky130_fd_sc_hd__clkbuf_2 hold1411 (.A(net2406),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[25] ),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(_2071_),
    .X(net2018));
 sky130_fd_sc_hd__buf_1 hold1414 (.A(net2408),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(_2034_),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(_2139_),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[11] ),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(_1972_),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[3] ),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[29] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[31] ),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(_2108_),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(_2109_),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(_2110_),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[28] ),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(_2088_),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(_2097_),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(_2098_),
    .X(net2032));
 sky130_fd_sc_hd__buf_1 hold1428 (.A(net2412),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(net109),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_0841_),
    .X(net748));
 sky130_fd_sc_hd__buf_2 hold1430 (.A(net2403),
    .X(net2035));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1431 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[15] ),
    .X(net2036));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1432 (.A(net2407),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[23] ),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(_1259_),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[17] ),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(_2009_),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(_2010_),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(_2012_),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(net124),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[8] ),
    .X(net749));
 sky130_fd_sc_hd__buf_2 hold1440 (.A(net2422),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(net100),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(net108),
    .X(net2047));
 sky130_fd_sc_hd__buf_2 hold1443 (.A(net2411),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(_3608_),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(_1369_),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(net120),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[10] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(_1961_),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(_1970_),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_0820_),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(_1971_),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(_1972_),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(net117),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(net122),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(net107),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[15] ),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(_1995_),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(_1996_),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(_1998_),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(net125),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[5] ),
    .X(net751));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1460 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[7] ),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[14] ),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(net111),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[4] ),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(net110),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(net118),
    .X(net2070));
 sky130_fd_sc_hd__buf_1 hold1466 (.A(net2413),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(net121),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(net126),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(net97),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0920_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(net105),
    .X(net2075));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1471 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[30] ),
    .X(net2076));
 sky130_fd_sc_hd__buf_2 hold1472 (.A(net2417),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(net106),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(net99),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(net113),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(net98),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(net112),
    .X(net2082));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1478 (.A(net2424),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(_3613_),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[9] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(_1374_),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(net104),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[1] ),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(net101),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(net103),
    .X(net2089));
 sky130_fd_sc_hd__buf_2 hold1485 (.A(net2430),
    .X(net2090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(_1368_),
    .X(net2091));
 sky130_fd_sc_hd__clkbuf_2 hold1487 (.A(net2106),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(net116),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(\U_DATAPATH.U_EX_MEM.o_rd_M[2] ),
    .X(net2094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_0821_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(_0915_),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(net115),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(net114),
    .X(net2097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(net119),
    .X(net2098));
 sky130_fd_sc_hd__buf_1 hold1494 (.A(net2421),
    .X(net2099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[4][2] ),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(_1080_),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[0] ),
    .X(net2102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(net123),
    .X(net2103));
 sky130_fd_sc_hd__buf_1 hold1499 (.A(net2418),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[17] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[27] ),
    .X(net755));
 sky130_fd_sc_hd__buf_1 hold1500 (.A(net2415),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[23] ),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(_0916_),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(net102),
    .X(net2108));
 sky130_fd_sc_hd__buf_2 hold1504 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[24] ),
    .X(net2109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(_3614_),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(\U_DATAPATH.U_EX_MEM.i_mem_write_EX ),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(_0913_),
    .X(net2112));
 sky130_fd_sc_hd__buf_1 hold1508 (.A(net2420),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(\U_CONTROL_UNIT.i_jump_EX ),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_0839_),
    .X(net756));
 sky130_fd_sc_hd__buf_4 hold1510 (.A(_1907_),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[29] ),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(net176),
    .X(net2117));
 sky130_fd_sc_hd__buf_1 hold1513 (.A(net2410),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[8][3] ),
    .X(net2119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(_1209_),
    .X(net2120));
 sky130_fd_sc_hd__buf_1 hold1516 (.A(net2414),
    .X(net2121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[2] ),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][1] ),
    .X(net2123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(_1301_),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[13] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[17] ),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(_0896_),
    .X(net2126));
 sky130_fd_sc_hd__clkbuf_4 hold1522 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[0] ),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(_3627_),
    .X(net2128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(_1387_),
    .X(net2129));
 sky130_fd_sc_hd__buf_1 hold1525 (.A(net2426),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(_1909_),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(_1911_),
    .X(net2132));
 sky130_fd_sc_hd__clkbuf_2 hold1528 (.A(net2402),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[1][0] ),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_0825_),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(_1268_),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[2] ),
    .X(net2136));
 sky130_fd_sc_hd__clkbuf_2 hold1532 (.A(net2401),
    .X(net2137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[24] ),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(_1481_),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[7] ),
    .X(net2140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(_1939_),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(_1949_),
    .X(net2142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(_1950_),
    .X(net2143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(_1951_),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[25] ),
    .X(net759));
 sky130_fd_sc_hd__buf_2 hold1540 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(_3625_),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(_1385_),
    .X(net2147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[29] ),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[31] ),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(_1582_),
    .X(net2150));
 sky130_fd_sc_hd__buf_1 hold1546 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[24] ),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(_2059_),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(_2060_),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(_2062_),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_0837_),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][17] ),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(_3571_),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(_1317_),
    .X(net2157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[14] ),
    .X(net2158));
 sky130_fd_sc_hd__buf_1 hold1554 (.A(_1804_),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[2] ),
    .X(net2160));
 sky130_fd_sc_hd__buf_1 hold1556 (.A(_1669_),
    .X(net2161));
 sky130_fd_sc_hd__clkbuf_2 hold1557 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[2] ),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[13] ),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(_1981_),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[1] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(_1990_),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(_1991_),
    .X(net2166));
 sky130_fd_sc_hd__clkbuf_2 hold1562 (.A(net2149),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[2][5] ),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(_1305_),
    .X(net2169));
 sky130_fd_sc_hd__buf_2 hold1565 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[3] ),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(_2702_),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1567 (.A(_3635_),
    .X(net2172));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1568 (.A(net2428),
    .X(net2173));
 sky130_fd_sc_hd__buf_1 hold1569 (.A(net2425),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_0948_),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_4 hold1570 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[28] ),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(_3610_),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[19] ),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(_2023_),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(_2024_),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(_2026_),
    .X(net2180));
 sky130_fd_sc_hd__clkbuf_4 hold1576 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[3] ),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(_3632_),
    .X(net2182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(_1396_),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[12] ),
    .X(net2184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[27] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(_1974_),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(_1983_),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(_1984_),
    .X(net2187));
 sky130_fd_sc_hd__clkbuf_4 hold1583 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[26] ),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(_3612_),
    .X(net2189));
 sky130_fd_sc_hd__clkbuf_2 hold1585 (.A(net2416),
    .X(net2190));
 sky130_fd_sc_hd__clkbuf_2 hold1586 (.A(net2404),
    .X(net2191));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1587 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[3] ),
    .X(net2192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(_1656_),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[27] ),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_0942_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(_2081_),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(_2082_),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(_2084_),
    .X(net2197));
 sky130_fd_sc_hd__buf_1 hold1593 (.A(net2427),
    .X(net2198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[16] ),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(_1508_),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[28] ),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(_2091_),
    .X(net2202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[3] ),
    .X(net2203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(_1917_),
    .X(net2204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0932_),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[30] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(_1921_),
    .X(net2205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[5] ),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(_1925_),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(_1926_),
    .X(net2208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(_1928_),
    .X(net2209));
 sky130_fd_sc_hd__buf_2 hold1605 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[1] ),
    .X(net2210));
 sky130_fd_sc_hd__clkbuf_2 hold1606 (.A(_2682_),
    .X(net2211));
 sky130_fd_sc_hd__buf_1 hold1607 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[16] ),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(_2002_),
    .X(net2213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(_2003_),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_0945_),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(_2005_),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[6] ),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(_1933_),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(_1941_),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(_1942_),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1615 (.A(_1943_),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[7] ),
    .X(net2221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(_1733_),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[26] ),
    .X(net2223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(_2075_),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[30] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(_2076_),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(_2077_),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[22] ),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(_2044_),
    .X(net2228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(_2045_),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(_2047_),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[9] ),
    .X(net2231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(_1954_),
    .X(net2232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(_1955_),
    .X(net2233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(_1957_),
    .X(net2234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_0977_),
    .X(net768));
 sky130_fd_sc_hd__buf_1 hold1630 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[18] ),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[9] ),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(_1791_),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[1] ),
    .X(net2238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(_3617_),
    .X(net2239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1635 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[13] ),
    .X(net2240));
 sky130_fd_sc_hd__buf_1 hold1636 (.A(_1836_),
    .X(net2241));
 sky130_fd_sc_hd__buf_2 hold1637 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[2] ),
    .X(net2242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(_3616_),
    .X(net2243));
 sky130_fd_sc_hd__buf_1 hold1639 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[6] ),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[11] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(_1935_),
    .X(net2245));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1641 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs2Addr_ID[0] ),
    .X(net2246));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1642 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[13] ),
    .X(net2247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(\U_CONTROL_UNIT.i_branch_EX ),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[29] ),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(_2095_),
    .X(net2250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(_2103_),
    .X(net2251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(_2104_),
    .X(net2252));
 sky130_fd_sc_hd__clkbuf_2 hold1648 (.A(net2423),
    .X(net2253));
 sky130_fd_sc_hd__clkbuf_2 hold1649 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[0] ),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_0958_),
    .X(net770));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1650 (.A(_2700_),
    .X(net2255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[10] ),
    .X(net2256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(_1756_),
    .X(net2257));
 sky130_fd_sc_hd__clkbuf_4 hold1653 (.A(\U_CONTROL_UNIT.U_OP_DECODER.i_op[2] ),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[27] ),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[21] ),
    .X(net2260));
 sky130_fd_sc_hd__buf_1 hold1656 (.A(_1642_),
    .X(net2261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[28] ),
    .X(net2262));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1658 (.A(_1568_),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[3] ),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[19] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[22] ),
    .X(net2265));
 sky130_fd_sc_hd__buf_1 hold1661 (.A(_1607_),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[11] ),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(_1780_),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[31] ),
    .X(net2269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[23] ),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(_2051_),
    .X(net2271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(_2052_),
    .X(net2272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(_2054_),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[12] ),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_0934_),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(_1811_),
    .X(net2275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[21] ),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(_2037_),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(_2038_),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(_2040_),
    .X(net2279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[30] ),
    .X(net2280));
 sky130_fd_sc_hd__buf_1 hold1676 (.A(_1559_),
    .X(net2281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[27] ),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[23] ),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[19] ),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[10] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(_1547_),
    .X(net2285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[10] ),
    .X(net2286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(_1964_),
    .X(net2287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[18] ),
    .X(net2288));
 sky130_fd_sc_hd__buf_1 hold1684 (.A(_1535_),
    .X(net2289));
 sky130_fd_sc_hd__buf_1 hold1685 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[15] ),
    .X(net2290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_3[2] ),
    .X(net2291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[25] ),
    .X(net2292));
 sky130_fd_sc_hd__buf_1 hold1688 (.A(_1461_),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[7] ),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_0957_),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[8] ),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(_1765_),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[4] ),
    .X(net2297));
 sky130_fd_sc_hd__buf_1 hold1693 (.A(_1719_),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[6] ),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(_1710_),
    .X(net2300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[21] ),
    .X(net2301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[15] ),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(_1825_),
    .X(net2303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[22] ),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[21] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[16] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[20] ),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[1] ),
    .X(net2306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(_1693_),
    .X(net2307));
 sky130_fd_sc_hd__clkbuf_2 hold1703 (.A(_0880_),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[25] ),
    .X(net2309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(_2066_),
    .X(net2310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(_2067_),
    .X(net2311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(_2069_),
    .X(net2312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[26] ),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[4] ),
    .X(net2314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_0931_),
    .X(net776));
 sky130_fd_sc_hd__buf_1 hold1710 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[11] ),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(_1968_),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[26] ),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[1] ),
    .X(net2319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[20] ),
    .X(net2320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1716 (.A(_2030_),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[17] ),
    .X(net2322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[29] ),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[5] ),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[16] ),
    .X(net777));
 sky130_fd_sc_hd__buf_1 hold1720 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[20] ),
    .X(net2325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(_2033_),
    .X(net2326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(\U_DATAPATH.U_ID_EX.o_rs2_EX[0] ),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[25] ),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[23] ),
    .X(net2329));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1725 (.A(\U_DATAPATH.U_ID_EX.o_alu_src_EX ),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(_1488_),
    .X(net2331));
 sky130_fd_sc_hd__clkbuf_2 hold1727 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[12] ),
    .X(net2332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(_1977_),
    .X(net2333));
 sky130_fd_sc_hd__clkbuf_4 hold1729 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[1] ),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_0828_),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[27] ),
    .X(net2335));
 sky130_fd_sc_hd__clkbuf_2 hold1731 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[3] ),
    .X(net2336));
 sky130_fd_sc_hd__clkbuf_2 hold1732 (.A(_2763_),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(_3058_),
    .X(net2338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(_0854_),
    .X(net2339));
 sky130_fd_sc_hd__clkbuf_2 hold1735 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[4] ),
    .X(net2340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(_1901_),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1737 (.A(_2780_),
    .X(net2342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(_0844_),
    .X(net2343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[8] ),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[29] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(_1772_),
    .X(net2345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(_0852_),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[29] ),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[16] ),
    .X(net2348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1744 (.A(_1513_),
    .X(net2349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1745 (.A(_0860_),
    .X(net2350));
 sky130_fd_sc_hd__buf_2 hold1746 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[2] ),
    .X(net2351));
 sky130_fd_sc_hd__clkbuf_4 hold1747 (.A(\U_DATAPATH.U_HAZARD_UNIT.i_rs1Addr_ID[0] ),
    .X(net2352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1748 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[31] ),
    .X(net2353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(_1596_),
    .X(net2354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_0976_),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1750 (.A(_0875_),
    .X(net2355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[9] ),
    .X(net2356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(_1795_),
    .X(net2357));
 sky130_fd_sc_hd__clkbuf_2 hold1753 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .X(net2358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(_0850_),
    .X(net2359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1755 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[18] ),
    .X(net2360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1756 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[20] ),
    .X(net2361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[28] ),
    .X(net2362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[26] ),
    .X(net2363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1759 (.A(_1471_),
    .X(net2364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[30] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1760 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[25] ),
    .X(net2365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1761 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[19] ),
    .X(net2366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1762 (.A(_1550_),
    .X(net2367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1763 (.A(_0863_),
    .X(net2368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1764 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[12] ),
    .X(net2369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1765 (.A(_1815_),
    .X(net2370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1766 (.A(_0856_),
    .X(net2371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1767 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[14] ),
    .X(net2372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1768 (.A(_1802_),
    .X(net2373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1769 (.A(_3134_),
    .X(net2374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_0842_),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1770 (.A(_0858_),
    .X(net2375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1771 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[21] ),
    .X(net2376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1772 (.A(_1640_),
    .X(net2377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1773 (.A(_0865_),
    .X(net2378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1774 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[2] ),
    .X(net2379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1775 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[7] ),
    .X(net2380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1776 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[13] ),
    .X(net2381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1777 (.A(_0857_),
    .X(net2382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1778 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[17] ),
    .X(net2383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1779 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[15] ),
    .X(net2384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[21] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1780 (.A(_1823_),
    .X(net2385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1781 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[30] ),
    .X(net2386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1782 (.A(_1562_),
    .X(net2387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1783 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[5] ),
    .X(net2388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1784 (.A(_1747_),
    .X(net2389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1785 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[23] ),
    .X(net2390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1786 (.A(_1629_),
    .X(net2391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1787 (.A(_0867_),
    .X(net2392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1788 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[22] ),
    .X(net2393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1789 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[1] ),
    .X(net2394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_0595_),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1790 (.A(_2824_),
    .X(net2395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1791 (.A(\U_DATAPATH.U_ID_EX.o_rs1_EX[4] ),
    .X(net2396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1792 (.A(\U_DATAPATH.U_ID_EX.o_imm_ex_EX[11] ),
    .X(net2397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1793 (.A(_1783_),
    .X(net2398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1794 (.A(\U_DATAPATH.U_EX_MEM.o_reg_write_M ),
    .X(net2399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1795 (.A(\U_DATAPATH.U_ID_EX.o_alu_ctrl_EX[2] ),
    .X(net2400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1796 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[12] ),
    .X(net2401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1797 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[8] ),
    .X(net2402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1798 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[27] ),
    .X(net2403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1799 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[9] ),
    .X(net2404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0833_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[13] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1800 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[17] ),
    .X(net2405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1801 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[24] ),
    .X(net2406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1802 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[22] ),
    .X(net2407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1803 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[20] ),
    .X(net2408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1804 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[1] ),
    .X(net2409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1805 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[3] ),
    .X(net2410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1806 (.A(\U_CONTROL_UNIT.U_ALU_DECODER.i_funct_7_5 ),
    .X(net2411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1807 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[10] ),
    .X(net2412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1808 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[11] ),
    .X(net2413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1809 (.A(\U_DATAPATH.U_ID_EX.i_rd_ID[2] ),
    .X(net2414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_0928_),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1810 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[25] ),
    .X(net2415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1811 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[26] ),
    .X(net2416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1812 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[29] ),
    .X(net2417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1813 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[16] ),
    .X(net2418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1814 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[27] ),
    .X(net2419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1815 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[19] ),
    .X(net2420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1816 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[21] ),
    .X(net2421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1817 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[20] ),
    .X(net2422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1818 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[28] ),
    .X(net2423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1819 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[25] ),
    .X(net2424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[0] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1820 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[15] ),
    .X(net2425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1821 (.A(\U_DATAPATH.U_ID_EX.o_pc_EX[2] ),
    .X(net2426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1822 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[11] ),
    .X(net2427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1823 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[4] ),
    .X(net2428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1824 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[19] ),
    .X(net2429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1825 (.A(\U_DATAPATH.U_IF_ID.o_instr_ID[31] ),
    .X(net2430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_0947_),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[4] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_0919_),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[31] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_0843_),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[27] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_0974_),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[19] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\U_DATAPATH.U_EX_MEM.i_reg_write_EX ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_0878_),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[6] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_0921_),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[3] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_0918_),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\U_DATAPATH.U_EX_MEM.o_result_src_M[0] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_0290_),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[22] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_0596_),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0922_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0966_),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[23] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_0835_),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[18] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_0830_),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[20] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_0594_),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[19] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_0831_),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[18] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_0622_),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[22] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[7] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_0819_),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[6] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_0326_),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[4] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_0608_),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[23] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_0597_),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[9] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_0613_),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0969_),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[21] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_0968_),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[5] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_0609_),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][0] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0778_),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][2] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_1144_),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][0] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_0540_),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[17] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][3] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_0479_),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[5] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_0325_),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[4] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_0578_),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[21] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_0936_),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][2] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_0510_),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0964_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][1] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_0747_),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][1] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_1175_),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[11] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_0585_),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][1] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_0541_),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[8] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_0612_),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[29] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[22] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_0626_),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][2] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_1112_),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][3] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_0447_),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\U_DATAPATH.U_EX_MEM.i_rd_EX[3] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_0813_),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][2] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_0542_),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0944_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][2] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_0748_),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][1] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_1143_),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][0] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(_0508_),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[27] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_0347_),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[3] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_0607_),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[22] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[7] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(_0611_),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[10] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_0584_),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][0] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_1110_),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][3] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(_0781_),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[7] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(_0581_),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0834_),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][3] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_1048_),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[2] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_0606_),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][3] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_0415_),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][2] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_0414_),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[26] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_0600_),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[25] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][3] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_0543_),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[8] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_0582_),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[13] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_0617_),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[24] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_0598_),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][0] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_1174_),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[6] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0940_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][1] ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(_0477_),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[25] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(_0629_),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][2] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(_1047_),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[24] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(_0628_),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[28] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_0602_),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[24] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[20] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(_0624_),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][0] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(_0746_),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[6] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(_0580_),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[16] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_0590_),
    .X(net922));
 sky130_fd_sc_hd__buf_1 hold318 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[2] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(_0091_),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0939_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[2] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(_0576_),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\U_DATAPATH.U_EX_MEM.i_pc_target_EX[1] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(_0715_),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[23] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(_0627_),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[12] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_0586_),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[30] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_0634_),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[26] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[5] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_0579_),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[12] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_0616_),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][0] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(_0444_),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[31] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(_0605_),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[13] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(_0587_),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0941_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[27] ),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(_0601_),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][12] ),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(_1122_),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][1] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(_0413_),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[17] ),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(_0591_),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\U_DATAPATH.U_EX_MEM.i_pc_target_EX[0] ),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(_0714_),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[4] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[29] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(_0603_),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][0] ),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(_0476_),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][26] ),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(_0804_),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[10] ),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(_0614_),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][1] ),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(_0445_),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0816_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][3] ),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(_0511_),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[14] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(_0618_),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[9] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(_0583_),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][8] ),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(_1118_),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[14] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(_0588_),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[15] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][10] ),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(_1120_),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][25] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(_0501_),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[16] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(_0620_),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][25] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(_0469_),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][20] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(_1194_),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0962_),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[18] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(_0592_),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[11] ),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(_0615_),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[30] ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(_0604_),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][25] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(_1070_),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[17] ),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(_0621_),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[15] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[15] ),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(_0619_),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][6] ),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(_0752_),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][20] ),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(_0464_),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][25] ),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(_0803_),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][11] ),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(_0519_),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0953_),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0930_),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][18] ),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(_0796_),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][16] ),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(_0556_),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][8] ),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(_1053_),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][12] ),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(_1186_),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[3] ),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(_0577_),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[26] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][29] ),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(_0537_),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_2 hold412 (.A(net2001),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][10] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_0518_),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][9] ),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_0549_),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][6] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_1116_),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][16] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0973_),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_0460_),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][8] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_0516_),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][24] ),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_0564_),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][6] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_1180_),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][10] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_1152_),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][21] ),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[21] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_0465_),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][12] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_0790_),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][4] ),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(_1178_),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][5] ),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_1147_),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][20] ),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_0798_),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][12] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0625_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_1154_),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][21] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_0561_),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][1] ),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_0779_),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][21] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_1195_),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][16] ),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_0428_),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][24] ),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[3] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_0468_),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][13] ),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_1123_),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][27] ),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(_0471_),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][27] ),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(_1072_),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][15] ),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(_0761_),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][14] ),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0950_),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_1124_),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][24] ),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(_1134_),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][1] ),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_0509_),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][20] ),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(_0766_),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][27] ),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(_0439_),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][1] ),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[25] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_1111_),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][21] ),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(_0529_),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][5] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(_0417_),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][20] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(_1130_),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][25] ),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(_1199_),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][30] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0972_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(_0474_),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][18] ),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(_0462_),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][2] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(_1176_),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][14] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(_1188_),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][31] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(_0539_),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][14] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[14] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_0458_),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][8] ),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_0786_),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[29] ),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_0633_),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][18] ),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(_0764_),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][21] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(_0799_),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[19] ),
    .X(net1104));
 sky130_fd_sc_hd__buf_1 hold5 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[3] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0826_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_0623_),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][26] ),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_0438_),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][5] ),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_0751_),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][15] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_0427_),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][26] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_0772_),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][16] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[28] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_1190_),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][15] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(_0523_),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][9] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(_0755_),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][23] ),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_0563_),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][10] ),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_0454_),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][30] ),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0840_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_0506_),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][20] ),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_0496_),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][16] ),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_0492_),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[6] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_0610_),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][23] ),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_1133_),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][3] ),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[23] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_1113_),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][30] ),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_0538_),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][10] ),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_0788_),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][23] ),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_0467_),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][23] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_1165_),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][23] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0970_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_0769_),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][5] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_0481_),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][0] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_0412_),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][9] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_0453_),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[15] ),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_0589_),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][26] ),
    .X(net1154));
 sky130_fd_sc_hd__buf_1 hold55 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[5] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_0470_),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][9] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_1151_),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][30] ),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_0570_),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][26] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_1168_),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][11] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_0551_),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][26] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0096_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_0566_),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][15] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_0555_),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][26] ),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_0502_),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][14] ),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_0792_),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][18] ),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_0558_),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][28] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[16] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_1138_),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][26] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_1136_),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][9] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_1119_),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][11] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_1185_),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][18] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_0494_),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][2] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0963_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_1338_),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][8] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_1150_),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][16] ),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_1158_),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][8] ),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_1182_),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][19] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_1129_),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][4] ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[24] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_0782_),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][7] ),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_1149_),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][16] ),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(_0524_),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][12] ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_0456_),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][10] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_0486_),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][23] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0094_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0971_),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_1197_),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][14] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_1156_),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][24] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_0436_),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][29] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(_0807_),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][15] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_0459_),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][23] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[28] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_0435_),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][12] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_0758_),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][28] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_0806_),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][25] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_0565_),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][31] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_1205_),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][10] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0943_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_1184_),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][11] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_0423_),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][6] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_0546_),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][18] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_1160_),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][18] ),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_0526_),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][15] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[27] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(_0491_),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][22] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(_1132_),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][31] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(_1076_),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][31] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(_1173_),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\U_DATAPATH.U_IF_ID.i_pcplus4_IF[14] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(_0334_),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][21] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0631_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_0433_),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][19] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(_0495_),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][17] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_1191_),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][29] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(_1074_),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][0] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(_1045_),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][11] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[26] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_0455_),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][8] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(_0754_),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][29] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_1171_),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][14] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_0760_),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][22] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(_1196_),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][6] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0630_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_0784_),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][23] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(_0801_),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][5] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(_1179_),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][12] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_0488_),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][6] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(_0418_),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][12] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[28] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(_0424_),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][31] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(_0809_),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][20] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_0432_),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][15] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(_1189_),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][22] ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(_0466_),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][24] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0632_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(_0500_),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][14] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(_1059_),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][21] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(_0767_),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][21] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(_1131_),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][7] ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(_1343_),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][31] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[12] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(_0777_),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][4] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(_1114_),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][22] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(_0530_),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][2] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(_0780_),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][6] ),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(_1342_),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][19] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[11] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0927_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(_0559_),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][28] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(_0472_),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][15] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(_1157_),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\U_DATAPATH.U_ID_EX.i_pc_ID[31] ),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(_0635_),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][16] ),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(_1126_),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][30] ),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[5] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(_0808_),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][31] ),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(_0571_),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][24] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(_0532_),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][3] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(_1145_),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[19] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(_0593_),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][10] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0952_),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(_1346_),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][4] ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(_1340_),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][1] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(_1046_),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][4] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(_0512_),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][4] ),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(_0750_),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][7] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[23] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(_1052_),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][8] ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(_1344_),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][9] ),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(_1183_),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][30] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(_0442_),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\U_DATAPATH.U_EX_MEM.i_result_src_EX[0] ),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(_0876_),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][19] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0938_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(_0765_),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][23] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(_1359_),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][14] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(_1350_),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][27] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(_0503_),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][28] ),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(_0504_),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][20] ),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[2] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(_0560_),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][14] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(_0426_),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][5] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(_0449_),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][30] ),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(_1172_),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][5] ),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(_1115_),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][25] ),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0917_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(_0437_),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][27] ),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(_0773_),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][22] ),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(_0800_),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][11] ),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(_0757_),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][0] ),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(_1142_),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][29] ),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[15] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(_0569_),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][28] ),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(_1170_),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][6] ),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(_1148_),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][2] ),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(_0446_),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][25] ),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(_0533_),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][16] ),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0827_),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(_0762_),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][8] ),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(_0484_),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][5] ),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(_0513_),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][10] ),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(_0756_),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][6] ),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(_0482_),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][28] ),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[26] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(_0568_),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][22] ),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(_0498_),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][22] ),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(_1164_),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][27] ),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(_1201_),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][24] ),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(_1166_),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][28] ),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0926_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0838_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(_1202_),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][6] ),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(_0450_),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][25] ),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(_1135_),
    .X(net1409));
 sky130_fd_sc_hd__buf_1 hold805 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[0] ),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(_0069_),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][17] ),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(_0557_),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][17] ),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[31] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(_0429_),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][21] ),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(_0497_),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][27] ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(_0567_),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][23] ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(_0499_),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][7] ),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(_1181_),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][15] ),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0978_),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(_0793_),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][9] ),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(_0421_),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][11] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(_0487_),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][5] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(_0783_),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][16] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(_1352_),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][16] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[9] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(_0794_),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][28] ),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(_0774_),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][18] ),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(_0430_),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][13] ),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(_0791_),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][10] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(_1055_),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][18] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0924_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(_1128_),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][31] ),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(_1141_),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][16] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(_1061_),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][13] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(_1187_),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][26] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(_1362_),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][22] ),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\U_DATAPATH.U_EX_MEM.i_pc_plus4_EX[10] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(_0434_),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][11] ),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(_1056_),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][18] ),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(_1192_),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][17] ),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(_1127_),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][10] ),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(_0422_),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][4] ),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0822_),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(_0448_),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][31] ),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(_0507_),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][11] ),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(_1153_),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][6] ),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(_0514_),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][11] ),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(_1121_),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][23] ),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[28] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(_1068_),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][24] ),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(_0802_),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][8] ),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(_0452_),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][14] ),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(_0554_),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][13] ),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(_1349_),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][25] ),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0975_),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(_0771_),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][19] ),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(_1193_),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[13] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(_0912_),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][17] ),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(_0763_),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][27] ),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(_0805_),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][19] ),
    .X(net1494));
 sky130_fd_sc_hd__buf_1 hold89 (.A(net2429),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(_0797_),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][3] ),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(_1177_),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][1] ),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(_1337_),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][29] ),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(_1365_),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][27] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(_0535_),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][10] ),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[13] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_3619_),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(_0550_),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][23] ),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(_0531_),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][30] ),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(_1366_),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][15] ),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(_1125_),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][14] ),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(_0522_),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][22] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_1380_),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(_1358_),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][11] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(_0789_),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][18] ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(_1354_),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][13] ),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(_0521_),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][31] ),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(_0443_),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][5] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\U_DATAPATH.U_EX_MEM.o_pc_plus4_M[20] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(_0545_),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][26] ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(_1071_),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][14] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(_0490_),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][7] ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(_1117_),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][17] ),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(_0461_),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][7] ),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0935_),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(_0753_),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][13] ),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(_0425_),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][26] ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(_1200_),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][25] ),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(_1361_),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][12] ),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(_1057_),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[3][24] ),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[9] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(_1198_),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][6] ),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(_1051_),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][21] ),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(_1066_),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][22] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(_0562_),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][30] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(_0776_),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][26] ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_0956_),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(_0534_),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][12] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(_1348_),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\U_DATAPATH.U_EX_MEM.o_alu_result_M[6] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(_0097_),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][28] ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(_0440_),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][19] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(_0527_),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][7] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\U_DATAPATH.U_EX_MEM.o_pc_target_M[12] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(_0547_),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[9][17] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(_0795_),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][30] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(_1075_),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][9] ),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(_0485_),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][31] ),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(_0475_),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][20] ),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0959_),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(_1162_),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[5][27] ),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(_1137_),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[6][27] ),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(_1169_),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][19] ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(_0463_),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[15][13] ),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(_0553_),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[10][13] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\U_DATAPATH.U_ID_EX.i_pc_plus4_ID[25] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(_0489_),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][17] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(_1062_),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][31] ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(_1367_),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][28] ),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(_0536_),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][18] ),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(_1063_),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[11][7] ),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0599_),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(_0451_),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[12][24] ),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(_1069_),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[0][15] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(_1351_),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[13][17] ),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(_0525_),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[14][19] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(_0431_),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\U_DATAPATH.U_STAGE_DECODE.U_REGISTER_FILE.registers[7][3] ),
    .X(net1604));
 sky130_fd_sc_hd__buf_1 input1 (.A(i_instr_ID[10]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(i_instr_ID[19]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(i_instr_ID[20]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(i_instr_ID[21]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(i_instr_ID[22]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(i_instr_ID[23]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(i_instr_ID[24]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(i_instr_ID[25]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(i_instr_ID[26]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(i_instr_ID[27]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(i_instr_ID[28]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(i_instr_ID[11]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(i_instr_ID[29]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(i_instr_ID[2]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(i_instr_ID[30]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(i_instr_ID[31]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(i_instr_ID[3]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(i_instr_ID[4]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input26 (.A(i_instr_ID[5]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(i_instr_ID[6]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(i_instr_ID[7]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(i_instr_ID[8]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input3 (.A(i_instr_ID[12]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(i_instr_ID[9]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(i_read_data_M[0]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(i_read_data_M[10]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(i_read_data_M[11]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(i_read_data_M[12]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(i_read_data_M[13]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(i_read_data_M[14]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(i_read_data_M[15]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(i_read_data_M[16]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(i_read_data_M[17]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input4 (.A(i_instr_ID[13]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(i_read_data_M[18]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(i_read_data_M[19]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(i_read_data_M[1]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(i_read_data_M[20]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(i_read_data_M[21]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(i_read_data_M[22]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(i_read_data_M[23]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(i_read_data_M[24]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(i_read_data_M[25]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(i_read_data_M[26]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(i_instr_ID[14]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(i_read_data_M[27]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(i_read_data_M[28]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(i_read_data_M[29]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(i_read_data_M[2]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(i_read_data_M[30]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(i_read_data_M[31]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(i_read_data_M[3]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(i_read_data_M[4]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(i_read_data_M[5]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(i_read_data_M[6]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(i_instr_ID[15]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(i_read_data_M[7]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(i_read_data_M[8]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(i_read_data_M[9]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_8 input63 (.A(rst),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input7 (.A(i_instr_ID[16]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(i_instr_ID[17]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(i_instr_ID[18]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 max_cap355 (.A(_2760_),
    .X(net355));
 sky130_fd_sc_hd__buf_12 output100 (.A(net100),
    .X(o_pc_IF[13]));
 sky130_fd_sc_hd__buf_12 output101 (.A(net101),
    .X(o_pc_IF[14]));
 sky130_fd_sc_hd__buf_12 output102 (.A(net102),
    .X(o_pc_IF[15]));
 sky130_fd_sc_hd__buf_12 output103 (.A(net103),
    .X(o_pc_IF[16]));
 sky130_fd_sc_hd__buf_12 output104 (.A(net104),
    .X(o_pc_IF[17]));
 sky130_fd_sc_hd__buf_12 output105 (.A(net105),
    .X(o_pc_IF[18]));
 sky130_fd_sc_hd__buf_12 output106 (.A(net106),
    .X(o_pc_IF[19]));
 sky130_fd_sc_hd__buf_12 output107 (.A(net107),
    .X(o_pc_IF[20]));
 sky130_fd_sc_hd__buf_12 output108 (.A(net108),
    .X(o_pc_IF[21]));
 sky130_fd_sc_hd__buf_12 output109 (.A(net109),
    .X(o_pc_IF[22]));
 sky130_fd_sc_hd__buf_12 output110 (.A(net110),
    .X(o_pc_IF[23]));
 sky130_fd_sc_hd__buf_12 output111 (.A(net111),
    .X(o_pc_IF[24]));
 sky130_fd_sc_hd__buf_12 output112 (.A(net112),
    .X(o_pc_IF[25]));
 sky130_fd_sc_hd__buf_12 output113 (.A(net113),
    .X(o_pc_IF[26]));
 sky130_fd_sc_hd__buf_12 output114 (.A(net114),
    .X(o_pc_IF[27]));
 sky130_fd_sc_hd__buf_12 output115 (.A(net115),
    .X(o_pc_IF[28]));
 sky130_fd_sc_hd__buf_12 output116 (.A(net116),
    .X(o_pc_IF[29]));
 sky130_fd_sc_hd__buf_12 output117 (.A(net117),
    .X(o_pc_IF[2]));
 sky130_fd_sc_hd__buf_12 output118 (.A(net118),
    .X(o_pc_IF[30]));
 sky130_fd_sc_hd__buf_12 output119 (.A(net119),
    .X(o_pc_IF[31]));
 sky130_fd_sc_hd__buf_12 output120 (.A(net120),
    .X(o_pc_IF[3]));
 sky130_fd_sc_hd__buf_12 output121 (.A(net121),
    .X(o_pc_IF[4]));
 sky130_fd_sc_hd__buf_12 output122 (.A(net122),
    .X(o_pc_IF[5]));
 sky130_fd_sc_hd__buf_12 output123 (.A(net123),
    .X(o_pc_IF[6]));
 sky130_fd_sc_hd__buf_12 output124 (.A(net124),
    .X(o_pc_IF[7]));
 sky130_fd_sc_hd__buf_12 output125 (.A(net125),
    .X(o_pc_IF[8]));
 sky130_fd_sc_hd__buf_12 output126 (.A(net126),
    .X(o_pc_IF[9]));
 sky130_fd_sc_hd__buf_12 output127 (.A(net127),
    .X(o_write_data_M[0]));
 sky130_fd_sc_hd__buf_12 output128 (.A(net128),
    .X(o_write_data_M[10]));
 sky130_fd_sc_hd__buf_12 output129 (.A(net129),
    .X(o_write_data_M[11]));
 sky130_fd_sc_hd__buf_12 output130 (.A(net130),
    .X(o_write_data_M[12]));
 sky130_fd_sc_hd__buf_12 output131 (.A(net131),
    .X(o_write_data_M[13]));
 sky130_fd_sc_hd__buf_12 output132 (.A(net132),
    .X(o_write_data_M[14]));
 sky130_fd_sc_hd__buf_12 output133 (.A(net133),
    .X(o_write_data_M[15]));
 sky130_fd_sc_hd__buf_12 output134 (.A(net134),
    .X(o_write_data_M[16]));
 sky130_fd_sc_hd__buf_12 output135 (.A(net135),
    .X(o_write_data_M[17]));
 sky130_fd_sc_hd__buf_12 output136 (.A(net136),
    .X(o_write_data_M[18]));
 sky130_fd_sc_hd__buf_12 output137 (.A(net137),
    .X(o_write_data_M[19]));
 sky130_fd_sc_hd__buf_12 output138 (.A(net138),
    .X(o_write_data_M[1]));
 sky130_fd_sc_hd__buf_12 output139 (.A(net139),
    .X(o_write_data_M[20]));
 sky130_fd_sc_hd__buf_12 output140 (.A(net140),
    .X(o_write_data_M[21]));
 sky130_fd_sc_hd__buf_12 output141 (.A(net141),
    .X(o_write_data_M[22]));
 sky130_fd_sc_hd__buf_12 output142 (.A(net142),
    .X(o_write_data_M[23]));
 sky130_fd_sc_hd__buf_12 output143 (.A(net143),
    .X(o_write_data_M[24]));
 sky130_fd_sc_hd__buf_12 output144 (.A(net144),
    .X(o_write_data_M[25]));
 sky130_fd_sc_hd__buf_12 output145 (.A(net145),
    .X(o_write_data_M[26]));
 sky130_fd_sc_hd__buf_12 output146 (.A(net146),
    .X(o_write_data_M[27]));
 sky130_fd_sc_hd__buf_12 output147 (.A(net147),
    .X(o_write_data_M[28]));
 sky130_fd_sc_hd__buf_12 output148 (.A(net148),
    .X(o_write_data_M[29]));
 sky130_fd_sc_hd__buf_12 output149 (.A(net149),
    .X(o_write_data_M[2]));
 sky130_fd_sc_hd__buf_12 output150 (.A(net150),
    .X(o_write_data_M[30]));
 sky130_fd_sc_hd__buf_12 output151 (.A(net151),
    .X(o_write_data_M[31]));
 sky130_fd_sc_hd__buf_12 output152 (.A(net152),
    .X(o_write_data_M[3]));
 sky130_fd_sc_hd__buf_12 output153 (.A(net153),
    .X(o_write_data_M[4]));
 sky130_fd_sc_hd__buf_12 output154 (.A(net154),
    .X(o_write_data_M[5]));
 sky130_fd_sc_hd__buf_12 output155 (.A(net155),
    .X(o_write_data_M[6]));
 sky130_fd_sc_hd__buf_12 output156 (.A(net156),
    .X(o_write_data_M[7]));
 sky130_fd_sc_hd__buf_12 output157 (.A(net157),
    .X(o_write_data_M[8]));
 sky130_fd_sc_hd__buf_12 output158 (.A(net158),
    .X(o_write_data_M[9]));
 sky130_fd_sc_hd__buf_12 output64 (.A(net64),
    .X(o_data_addr_M[0]));
 sky130_fd_sc_hd__buf_12 output65 (.A(net65),
    .X(o_data_addr_M[10]));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(o_data_addr_M[11]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(o_data_addr_M[12]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(o_data_addr_M[13]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(o_data_addr_M[14]));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(o_data_addr_M[15]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(o_data_addr_M[16]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net72),
    .X(o_data_addr_M[17]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(o_data_addr_M[18]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(o_data_addr_M[19]));
 sky130_fd_sc_hd__buf_12 output75 (.A(net75),
    .X(o_data_addr_M[1]));
 sky130_fd_sc_hd__buf_12 output76 (.A(net76),
    .X(o_data_addr_M[20]));
 sky130_fd_sc_hd__buf_12 output77 (.A(net77),
    .X(o_data_addr_M[21]));
 sky130_fd_sc_hd__buf_12 output78 (.A(net78),
    .X(o_data_addr_M[22]));
 sky130_fd_sc_hd__buf_12 output79 (.A(net79),
    .X(o_data_addr_M[23]));
 sky130_fd_sc_hd__buf_12 output80 (.A(net80),
    .X(o_data_addr_M[24]));
 sky130_fd_sc_hd__buf_12 output81 (.A(net81),
    .X(o_data_addr_M[25]));
 sky130_fd_sc_hd__buf_12 output82 (.A(net82),
    .X(o_data_addr_M[26]));
 sky130_fd_sc_hd__buf_12 output83 (.A(net83),
    .X(o_data_addr_M[27]));
 sky130_fd_sc_hd__buf_12 output84 (.A(net84),
    .X(o_data_addr_M[28]));
 sky130_fd_sc_hd__buf_12 output85 (.A(net85),
    .X(o_data_addr_M[29]));
 sky130_fd_sc_hd__buf_12 output86 (.A(net86),
    .X(o_data_addr_M[2]));
 sky130_fd_sc_hd__buf_12 output87 (.A(net87),
    .X(o_data_addr_M[30]));
 sky130_fd_sc_hd__buf_12 output88 (.A(net88),
    .X(o_data_addr_M[31]));
 sky130_fd_sc_hd__buf_12 output89 (.A(net89),
    .X(o_data_addr_M[3]));
 sky130_fd_sc_hd__buf_12 output90 (.A(net90),
    .X(o_data_addr_M[4]));
 sky130_fd_sc_hd__buf_12 output91 (.A(net91),
    .X(o_data_addr_M[5]));
 sky130_fd_sc_hd__buf_12 output92 (.A(net92),
    .X(o_data_addr_M[6]));
 sky130_fd_sc_hd__buf_12 output93 (.A(net93),
    .X(o_data_addr_M[7]));
 sky130_fd_sc_hd__buf_12 output94 (.A(net94),
    .X(o_data_addr_M[8]));
 sky130_fd_sc_hd__buf_12 output95 (.A(net95),
    .X(o_data_addr_M[9]));
 sky130_fd_sc_hd__buf_12 output96 (.A(net96),
    .X(o_mem_write_M));
 sky130_fd_sc_hd__buf_12 output97 (.A(net97),
    .X(o_pc_IF[10]));
 sky130_fd_sc_hd__buf_12 output98 (.A(net98),
    .X(o_pc_IF[11]));
 sky130_fd_sc_hd__buf_12 output99 (.A(net99),
    .X(o_pc_IF[12]));
 assign o_pc_IF[0] = net473;
 assign o_pc_IF[1] = net474;
endmodule

