// This is the unpowered netlist.
module uart_wbs_bridge (clk,
    i_start_rx,
    i_uart_rx,
    o_uart_tx,
    rst,
    wb_ack_i,
    wb_cyc_o,
    wb_stb_o,
    wb_we_o,
    wb_adr_o,
    wb_dat_i,
    wb_dat_o);
 input clk;
 input i_start_rx;
 input i_uart_rx;
 output o_uart_tx;
 input rst;
 input wb_ack_i;
 output wb_cyc_o;
 output wb_stb_o;
 output wb_we_o;
 output [15:0] wb_adr_o;
 input [31:0] wb_dat_i;
 output [31:0] wb_dat_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire \addr_reg[0] ;
 wire \addr_reg[10] ;
 wire \addr_reg[11] ;
 wire \addr_reg[12] ;
 wire \addr_reg[13] ;
 wire \addr_reg[14] ;
 wire \addr_reg[15] ;
 wire \addr_reg[1] ;
 wire \addr_reg[2] ;
 wire \addr_reg[3] ;
 wire \addr_reg[4] ;
 wire \addr_reg[5] ;
 wire \addr_reg[6] ;
 wire \addr_reg[7] ;
 wire \addr_reg[8] ;
 wire \addr_reg[9] ;
 wire \byte_count[0] ;
 wire \byte_count[1] ;
 wire \byte_count[2] ;
 wire \byte_count[3] ;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire \cmd_reg[0] ;
 wire \cmd_reg[1] ;
 wire \cmd_reg[2] ;
 wire \cmd_reg[3] ;
 wire \cmd_reg[4] ;
 wire \cmd_reg[5] ;
 wire \cmd_reg[6] ;
 wire \cmd_reg[7] ;
 wire \data_reg[0] ;
 wire \data_reg[10] ;
 wire \data_reg[11] ;
 wire \data_reg[12] ;
 wire \data_reg[13] ;
 wire \data_reg[14] ;
 wire \data_reg[15] ;
 wire \data_reg[16] ;
 wire \data_reg[17] ;
 wire \data_reg[18] ;
 wire \data_reg[19] ;
 wire \data_reg[1] ;
 wire \data_reg[20] ;
 wire \data_reg[21] ;
 wire \data_reg[22] ;
 wire \data_reg[23] ;
 wire \data_reg[2] ;
 wire \data_reg[3] ;
 wire \data_reg[4] ;
 wire \data_reg[5] ;
 wire \data_reg[6] ;
 wire \data_reg[7] ;
 wire \data_reg[8] ;
 wire \data_reg[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \uart_rx_inst.bit_index[0] ;
 wire \uart_rx_inst.bit_index[1] ;
 wire \uart_rx_inst.bit_index[2] ;
 wire \uart_rx_inst.bit_index[3] ;
 wire \uart_rx_inst.clock_count[0] ;
 wire \uart_rx_inst.clock_count[10] ;
 wire \uart_rx_inst.clock_count[11] ;
 wire \uart_rx_inst.clock_count[12] ;
 wire \uart_rx_inst.clock_count[13] ;
 wire \uart_rx_inst.clock_count[14] ;
 wire \uart_rx_inst.clock_count[15] ;
 wire \uart_rx_inst.clock_count[1] ;
 wire \uart_rx_inst.clock_count[2] ;
 wire \uart_rx_inst.clock_count[3] ;
 wire \uart_rx_inst.clock_count[4] ;
 wire \uart_rx_inst.clock_count[5] ;
 wire \uart_rx_inst.clock_count[6] ;
 wire \uart_rx_inst.clock_count[7] ;
 wire \uart_rx_inst.clock_count[8] ;
 wire \uart_rx_inst.clock_count[9] ;
 wire \uart_rx_inst.o_data[0] ;
 wire \uart_rx_inst.o_data[1] ;
 wire \uart_rx_inst.o_data[2] ;
 wire \uart_rx_inst.o_data[3] ;
 wire \uart_rx_inst.o_data[4] ;
 wire \uart_rx_inst.o_data[5] ;
 wire \uart_rx_inst.o_data[6] ;
 wire \uart_rx_inst.o_data[7] ;
 wire \uart_rx_inst.o_data_valid ;
 wire \uart_rx_inst.receiving ;
 wire \uart_rx_inst.rx_sync_1 ;
 wire \uart_rx_inst.rx_sync_2 ;
 wire \uart_rx_inst.shift_reg[0] ;
 wire \uart_rx_inst.shift_reg[1] ;
 wire \uart_rx_inst.shift_reg[2] ;
 wire \uart_rx_inst.shift_reg[3] ;
 wire \uart_rx_inst.shift_reg[4] ;
 wire \uart_rx_inst.shift_reg[5] ;
 wire \uart_rx_inst.shift_reg[6] ;
 wire \uart_rx_inst.shift_reg[7] ;
 wire \uart_tx_inst.bit_index[0] ;
 wire \uart_tx_inst.bit_index[1] ;
 wire \uart_tx_inst.bit_index[2] ;
 wire \uart_tx_inst.bit_index[3] ;
 wire \uart_tx_inst.clock_count[0] ;
 wire \uart_tx_inst.clock_count[10] ;
 wire \uart_tx_inst.clock_count[11] ;
 wire \uart_tx_inst.clock_count[12] ;
 wire \uart_tx_inst.clock_count[13] ;
 wire \uart_tx_inst.clock_count[14] ;
 wire \uart_tx_inst.clock_count[15] ;
 wire \uart_tx_inst.clock_count[1] ;
 wire \uart_tx_inst.clock_count[2] ;
 wire \uart_tx_inst.clock_count[3] ;
 wire \uart_tx_inst.clock_count[4] ;
 wire \uart_tx_inst.clock_count[5] ;
 wire \uart_tx_inst.clock_count[6] ;
 wire \uart_tx_inst.clock_count[7] ;
 wire \uart_tx_inst.clock_count[8] ;
 wire \uart_tx_inst.clock_count[9] ;
 wire \uart_tx_inst.i_data[0] ;
 wire \uart_tx_inst.i_data[1] ;
 wire \uart_tx_inst.i_data[2] ;
 wire \uart_tx_inst.i_data[3] ;
 wire \uart_tx_inst.i_data[4] ;
 wire \uart_tx_inst.i_data[5] ;
 wire \uart_tx_inst.i_data[6] ;
 wire \uart_tx_inst.i_data[7] ;
 wire \uart_tx_inst.i_data_valid ;
 wire \uart_tx_inst.o_ready ;
 wire \uart_tx_inst.shift_reg[1] ;
 wire \uart_tx_inst.shift_reg[2] ;
 wire \uart_tx_inst.shift_reg[3] ;
 wire \uart_tx_inst.shift_reg[4] ;
 wire \uart_tx_inst.shift_reg[5] ;
 wire \uart_tx_inst.shift_reg[6] ;
 wire \uart_tx_inst.shift_reg[7] ;
 wire \uart_tx_inst.shift_reg[8] ;
 wire \uart_tx_inst.shift_reg[9] ;
 wire \uart_tx_inst.transmitting ;

 sky130_fd_sc_hd__diode_2 ANTENNA__0618__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__B1 (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__B (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__A (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0724__A (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0739__A (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__B (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__S (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0756__S (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__S (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__S (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__S (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0760__S (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0761__S (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0762__S (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0766__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__A1 (.DIODE(\uart_rx_inst.o_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__A1 (.DIODE(\uart_rx_inst.o_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0770__A1 (.DIODE(\uart_rx_inst.o_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__A1 (.DIODE(\uart_rx_inst.o_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0831__C (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0841__D_N (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0862__A (.DIODE(\uart_rx_inst.o_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0862__B (.DIODE(\uart_rx_inst.o_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0862__D_N (.DIODE(\uart_rx_inst.o_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__A_N (.DIODE(\uart_rx_inst.o_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__C (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__D (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__0876__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0883__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0887__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0890__C_N (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0893__A1_N (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0893__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0895__A1_N (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__C_N (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__0897__A1_N (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0897__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0898__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0898__C_N (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__0899__A1_N (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0899__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0900__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0901__A1_N (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0901__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0902__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0902__C_N (.DIODE(\uart_rx_inst.o_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0903__A1_N (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0903__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0904__C_N (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__0905__A1_N (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0905__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0906__C_N (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__0907__A1_N (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0907__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0908__B (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0909__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0909__B1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0909__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__B1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__B2 (.DIODE(\uart_rx_inst.o_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0911__B1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0911__B2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__0912__B1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0912__B2 (.DIODE(\uart_rx_inst.o_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0913__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0913__B1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0913__B2 (.DIODE(\uart_rx_inst.o_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0914__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0914__B1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0914__B2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__B1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__0916__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0916__B1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0916__B2 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__B2 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0920__B2 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0922__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0922__B2 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0924__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0924__B2 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__B2 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0928__B2 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0932__B2 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0934__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0934__B1 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0934__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__0935__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0935__B1 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0935__B2 (.DIODE(\uart_rx_inst.o_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0936__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0936__B1 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0937__B1 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0937__B2 (.DIODE(\uart_rx_inst.o_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__B1 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__B2 (.DIODE(\uart_rx_inst.o_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0939__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0939__B1 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0939__B2 (.DIODE(\uart_rx_inst.o_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0940__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0940__B1 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0941__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0941__B1 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0941__B2 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__0943__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0944__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0946__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0947__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0948__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0950__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__0952__A0 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__0953__A0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__0955__A0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__0956__A0 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__0957__A0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__0960__S0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0960__S1 (.DIODE(\byte_count[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__S0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__S1 (.DIODE(\byte_count[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__S0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__S1 (.DIODE(\byte_count[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0969__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__0969__S0 (.DIODE(\byte_count[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0969__S1 (.DIODE(\byte_count[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0972__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__0972__S0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0972__S1 (.DIODE(\byte_count[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__S0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__S1 (.DIODE(\byte_count[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__A0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__S0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__S1 (.DIODE(\byte_count[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__S0 (.DIODE(\byte_count[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__S1 (.DIODE(\byte_count[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__B (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0989__B (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0993__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__0993__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0997__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__0997__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1002__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1003__S (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1005__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1006__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1007__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1011__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1013__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1014__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1017__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1018__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1019__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1020__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__A2 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1026__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1027__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1028__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1029__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1034__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1036__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1040__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1041__S (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1197__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1420__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold161_A (.DIODE(\byte_count[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold163_A (.DIODE(\uart_rx_inst.o_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold167_A (.DIODE(\uart_rx_inst.o_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold172_A (.DIODE(\uart_rx_inst.o_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold174_A (.DIODE(\uart_rx_inst.o_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold208_A (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold228_A (.DIODE(\byte_count[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold303_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold91_A (.DIODE(\byte_count[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net54));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__inv_2 _0617_ (.A(net400),
    .Y(_0372_));
 sky130_fd_sc_hd__inv_2 _0618_ (.A(net179),
    .Y(_0373_));
 sky130_fd_sc_hd__inv_2 _0619_ (.A(net225),
    .Y(_0374_));
 sky130_fd_sc_hd__inv_2 _0620_ (.A(net343),
    .Y(_0375_));
 sky130_fd_sc_hd__inv_2 _0621_ (.A(net171),
    .Y(_0376_));
 sky130_fd_sc_hd__inv_2 _0622_ (.A(net350),
    .Y(_0377_));
 sky130_fd_sc_hd__inv_2 _0623_ (.A(net412),
    .Y(_0378_));
 sky130_fd_sc_hd__inv_2 _0624_ (.A(net299),
    .Y(_0379_));
 sky130_fd_sc_hd__inv_2 _0625_ (.A(net256),
    .Y(_0380_));
 sky130_fd_sc_hd__inv_2 _0626_ (.A(net275),
    .Y(_0381_));
 sky130_fd_sc_hd__inv_2 _0627_ (.A(net4),
    .Y(_0382_));
 sky130_fd_sc_hd__inv_2 _0628_ (.A(net104),
    .Y(_0003_));
 sky130_fd_sc_hd__nor2_1 _0629_ (.A(net343),
    .B(net171),
    .Y(_0383_));
 sky130_fd_sc_hd__or2_2 _0630_ (.A(net343),
    .B(net171),
    .X(_0384_));
 sky130_fd_sc_hd__or2_2 _0631_ (.A(net193),
    .B(net225),
    .X(_0385_));
 sky130_fd_sc_hd__nor2_1 _0632_ (.A(_0384_),
    .B(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__o21a_1 _0633_ (.A1(net225),
    .A2(_0384_),
    .B1(net193),
    .X(_0387_));
 sky130_fd_sc_hd__or4bb_1 _0634_ (.A(net324),
    .B(net313),
    .C_N(net357),
    .D_N(net372),
    .X(_0388_));
 sky130_fd_sc_hd__or4bb_1 _0635_ (.A(net350),
    .B(net345),
    .C_N(net347),
    .D_N(\uart_rx_inst.clock_count[0] ),
    .X(_0389_));
 sky130_fd_sc_hd__or4b_1 _0636_ (.A(net309),
    .B(net412),
    .C(net328),
    .D_N(\uart_rx_inst.clock_count[6] ),
    .X(_0390_));
 sky130_fd_sc_hd__or4bb_1 _0637_ (.A(net336),
    .B(net326),
    .C_N(net340),
    .D_N(net380),
    .X(_0391_));
 sky130_fd_sc_hd__nor4_1 _0638_ (.A(_0388_),
    .B(net351),
    .C(net413),
    .D(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__nand2_2 _0639_ (.A(net97),
    .B(net95),
    .Y(_0393_));
 sky130_fd_sc_hd__nor2_1 _0640_ (.A(_0387_),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__or4bb_1 _0641_ (.A(_0386_),
    .B(_0387_),
    .C_N(net95),
    .D_N(net97),
    .X(_0395_));
 sky130_fd_sc_hd__or4_1 _0642_ (.A(_0388_),
    .B(_0389_),
    .C(_0390_),
    .D(_0391_),
    .X(_0396_));
 sky130_fd_sc_hd__or4b_4 _0643_ (.A(_0386_),
    .B(_0387_),
    .C(net352),
    .D_N(net97),
    .X(_0397_));
 sky130_fd_sc_hd__o31a_1 _0644_ (.A1(net225),
    .A2(_0384_),
    .A3(net353),
    .B1(net181),
    .X(_0398_));
 sky130_fd_sc_hd__nor2_1 _0645_ (.A(net343),
    .B(_0376_),
    .Y(_0399_));
 sky130_fd_sc_hd__xnor2_1 _0646_ (.A(net225),
    .B(net343),
    .Y(_0400_));
 sky130_fd_sc_hd__xor2_1 _0647_ (.A(net225),
    .B(net343),
    .X(_0401_));
 sky130_fd_sc_hd__o21a_1 _0648_ (.A1(_0384_),
    .A2(_0385_),
    .B1(net162),
    .X(_0402_));
 sky130_fd_sc_hd__nor2_1 _0649_ (.A(_0397_),
    .B(_0401_),
    .Y(_0403_));
 sky130_fd_sc_hd__a31o_1 _0650_ (.A1(_0383_),
    .A2(net163),
    .A3(_0403_),
    .B1(_0398_),
    .X(_0369_));
 sky130_fd_sc_hd__nor2_1 _0651_ (.A(_0375_),
    .B(_0376_),
    .Y(_0404_));
 sky130_fd_sc_hd__nand2_1 _0652_ (.A(net343),
    .B(net171),
    .Y(_0405_));
 sky130_fd_sc_hd__or2_1 _0653_ (.A(_0374_),
    .B(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__or2_1 _0654_ (.A(_0395_),
    .B(net226),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _0655_ (.A0(net162),
    .A1(net144),
    .S(_0407_),
    .X(_0368_));
 sky130_fd_sc_hd__nor2_1 _0656_ (.A(_0375_),
    .B(net171),
    .Y(_0408_));
 sky130_fd_sc_hd__or3b_1 _0657_ (.A(_0395_),
    .B(_0401_),
    .C_N(net172),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _0658_ (.A0(net162),
    .A1(net150),
    .S(net173),
    .X(_0367_));
 sky130_fd_sc_hd__o41a_1 _0659_ (.A1(_0374_),
    .A2(net343),
    .A3(_0376_),
    .A4(_0395_),
    .B1(net222),
    .X(_0410_));
 sky130_fd_sc_hd__a41o_1 _0660_ (.A1(net162),
    .A2(_0385_),
    .A3(_0394_),
    .A4(_0399_),
    .B1(_0410_),
    .X(_0366_));
 sky130_fd_sc_hd__o31a_1 _0661_ (.A1(_0374_),
    .A2(_0384_),
    .A3(net353),
    .B1(net266),
    .X(_0411_));
 sky130_fd_sc_hd__nor2_1 _0662_ (.A(_0397_),
    .B(_0400_),
    .Y(_0412_));
 sky130_fd_sc_hd__a31o_1 _0663_ (.A1(net162),
    .A2(_0383_),
    .A3(_0412_),
    .B1(_0411_),
    .X(_0365_));
 sky130_fd_sc_hd__o31a_1 _0664_ (.A1(_0385_),
    .A2(_0397_),
    .A3(_0405_),
    .B1(net183),
    .X(_0413_));
 sky130_fd_sc_hd__a31o_1 _0665_ (.A1(net162),
    .A2(_0404_),
    .A3(_0412_),
    .B1(_0413_),
    .X(_0364_));
 sky130_fd_sc_hd__o41a_1 _0666_ (.A1(_0375_),
    .A2(net171),
    .A3(_0397_),
    .A4(_0400_),
    .B1(net132),
    .X(_0414_));
 sky130_fd_sc_hd__a31o_1 _0667_ (.A1(net162),
    .A2(net172),
    .A3(_0412_),
    .B1(net354),
    .X(_0363_));
 sky130_fd_sc_hd__or3b_1 _0668_ (.A(_0385_),
    .B(_0397_),
    .C_N(_0399_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _0669_ (.A0(net163),
    .A1(net148),
    .S(_0415_),
    .X(_0362_));
 sky130_fd_sc_hd__nand2_1 _0670_ (.A(net384),
    .B(\uart_tx_inst.bit_index[0] ),
    .Y(_0416_));
 sky130_fd_sc_hd__and3_1 _0671_ (.A(net377),
    .B(net384),
    .C(\uart_tx_inst.bit_index[0] ),
    .X(_0417_));
 sky130_fd_sc_hd__or4bb_1 _0672_ (.A(net404),
    .B(net400),
    .C_N(net366),
    .D_N(net331),
    .X(_0418_));
 sky130_fd_sc_hd__or4bb_1 _0673_ (.A(net302),
    .B(net333),
    .C_N(net382),
    .D_N(net394),
    .X(_0419_));
 sky130_fd_sc_hd__or4b_1 _0674_ (.A(net396),
    .B(net402),
    .C(net391),
    .D_N(net359),
    .X(_0420_));
 sky130_fd_sc_hd__or4bb_1 _0675_ (.A(net407),
    .B(net315),
    .C_N(net362),
    .D_N(net368),
    .X(_0421_));
 sky130_fd_sc_hd__nor4_1 _0676_ (.A(_0418_),
    .B(_0419_),
    .C(_0420_),
    .D(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__nand2_1 _0677_ (.A(net96),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__and3_1 _0678_ (.A(net96),
    .B(_0417_),
    .C(_0422_),
    .X(_0424_));
 sky130_fd_sc_hd__nand2_2 _0679_ (.A(net386),
    .B(net410),
    .Y(_0425_));
 sky130_fd_sc_hd__a21oi_4 _0680_ (.A1(net386),
    .A2(net410),
    .B1(net96),
    .Y(_0426_));
 sky130_fd_sc_hd__or4_1 _0681_ (.A(_0418_),
    .B(_0419_),
    .C(_0420_),
    .D(_0421_),
    .X(_0427_));
 sky130_fd_sc_hd__and2_1 _0682_ (.A(net96),
    .B(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__a21oi_1 _0683_ (.A1(net96),
    .A2(_0427_),
    .B1(_0426_),
    .Y(_0429_));
 sky130_fd_sc_hd__or2_1 _0684_ (.A(_0426_),
    .B(_0428_),
    .X(_0430_));
 sky130_fd_sc_hd__o21ai_1 _0685_ (.A1(_0417_),
    .A2(_0423_),
    .B1(_0429_),
    .Y(_0431_));
 sky130_fd_sc_hd__mux2_1 _0686_ (.A0(_0424_),
    .A1(_0431_),
    .S(net388),
    .X(_0361_));
 sky130_fd_sc_hd__or3_1 _0687_ (.A(net377),
    .B(_0416_),
    .C(_0423_),
    .X(_0432_));
 sky130_fd_sc_hd__a21bo_1 _0688_ (.A1(net377),
    .A2(_0431_),
    .B1_N(_0432_),
    .X(_0360_));
 sky130_fd_sc_hd__or2_1 _0689_ (.A(net384),
    .B(\uart_tx_inst.bit_index[0] ),
    .X(_0433_));
 sky130_fd_sc_hd__nand2_1 _0690_ (.A(_0416_),
    .B(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__a2bb2o_1 _0691_ (.A1_N(_0423_),
    .A2_N(_0434_),
    .B1(_0430_),
    .B2(net384),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _0692_ (.A0(_0429_),
    .A1(_0423_),
    .S(net416),
    .X(_0358_));
 sky130_fd_sc_hd__and4_2 _0693_ (.A(net315),
    .B(net362),
    .C(net382),
    .D(net394),
    .X(_0435_));
 sky130_fd_sc_hd__inv_2 _0694_ (.A(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__nand2_1 _0695_ (.A(net368),
    .B(_0435_),
    .Y(_0437_));
 sky130_fd_sc_hd__and2_1 _0696_ (.A(net407),
    .B(net368),
    .X(_0438_));
 sky130_fd_sc_hd__and2_1 _0697_ (.A(_0435_),
    .B(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__and2_1 _0698_ (.A(net391),
    .B(net359),
    .X(_0440_));
 sky130_fd_sc_hd__and3_1 _0699_ (.A(_0435_),
    .B(_0438_),
    .C(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__and4_1 _0700_ (.A(net400),
    .B(net366),
    .C(net396),
    .D(\uart_tx_inst.clock_count[8] ),
    .X(_0442_));
 sky130_fd_sc_hd__and3_1 _0701_ (.A(net331),
    .B(_0441_),
    .C(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__and4_1 _0702_ (.A(\uart_tx_inst.clock_count[14] ),
    .B(\uart_tx_inst.clock_count[13] ),
    .C(net96),
    .D(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__nor2_8 _0703_ (.A(net96),
    .B(_0425_),
    .Y(_0445_));
 sky130_fd_sc_hd__or2_1 _0704_ (.A(net96),
    .B(_0425_),
    .X(_0446_));
 sky130_fd_sc_hd__a41oi_2 _0705_ (.A1(net333),
    .A2(\uart_tx_inst.clock_count[13] ),
    .A3(net96),
    .A4(_0443_),
    .B1(_0445_),
    .Y(_0447_));
 sky130_fd_sc_hd__and3_1 _0706_ (.A(net404),
    .B(net96),
    .C(_0443_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _0707_ (.A0(_0444_),
    .A1(_0447_),
    .S(net302),
    .X(_0357_));
 sky130_fd_sc_hd__o21a_1 _0708_ (.A1(net333),
    .A2(_0448_),
    .B1(_0447_),
    .X(_0356_));
 sky130_fd_sc_hd__a22oi_1 _0709_ (.A1(net96),
    .A2(_0443_),
    .B1(_0446_),
    .B2(net404),
    .Y(_0449_));
 sky130_fd_sc_hd__nor2_1 _0710_ (.A(_0448_),
    .B(net405),
    .Y(_0355_));
 sky130_fd_sc_hd__a21oi_1 _0711_ (.A1(_0441_),
    .A2(_0442_),
    .B1(net331),
    .Y(_0450_));
 sky130_fd_sc_hd__nor2_1 _0712_ (.A(_0443_),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__a22o_1 _0713_ (.A1(net331),
    .A2(_0426_),
    .B1(_0428_),
    .B2(_0451_),
    .X(_0354_));
 sky130_fd_sc_hd__and4_1 _0714_ (.A(net96),
    .B(_0435_),
    .C(_0438_),
    .D(_0440_),
    .X(_0452_));
 sky130_fd_sc_hd__and3_1 _0715_ (.A(net396),
    .B(\uart_tx_inst.clock_count[8] ),
    .C(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__nand2_1 _0716_ (.A(net366),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__nor2_1 _0717_ (.A(_0372_),
    .B(_0445_),
    .Y(_0455_));
 sky130_fd_sc_hd__mux2_1 _0718_ (.A0(_0372_),
    .A1(_0455_),
    .S(_0454_),
    .X(_0353_));
 sky130_fd_sc_hd__and4b_1 _0719_ (.A_N(_0426_),
    .B(_0441_),
    .C(\uart_tx_inst.clock_count[9] ),
    .D(\uart_tx_inst.clock_count[8] ),
    .X(_0456_));
 sky130_fd_sc_hd__nor2_1 _0720_ (.A(_0429_),
    .B(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__mux2_1 _0721_ (.A0(_0453_),
    .A1(_0457_),
    .S(net366),
    .X(_0352_));
 sky130_fd_sc_hd__a21oi_1 _0722_ (.A1(\uart_tx_inst.clock_count[8] ),
    .A2(_0452_),
    .B1(net396),
    .Y(_0458_));
 sky130_fd_sc_hd__nor3_1 _0723_ (.A(_0445_),
    .B(_0453_),
    .C(net397),
    .Y(_0351_));
 sky130_fd_sc_hd__nor2_1 _0724_ (.A(_0445_),
    .B(_0452_),
    .Y(_0459_));
 sky130_fd_sc_hd__mux2_1 _0725_ (.A0(_0452_),
    .A1(_0459_),
    .S(net402),
    .X(_0350_));
 sky130_fd_sc_hd__nand2_1 _0726_ (.A(net96),
    .B(_0439_),
    .Y(_0460_));
 sky130_fd_sc_hd__a31o_1 _0727_ (.A1(net359),
    .A2(net96),
    .A3(_0439_),
    .B1(net391),
    .X(_0461_));
 sky130_fd_sc_hd__and2_1 _0728_ (.A(_0459_),
    .B(net392),
    .X(_0349_));
 sky130_fd_sc_hd__nand2b_1 _0729_ (.A_N(_0426_),
    .B(_0439_),
    .Y(_0462_));
 sky130_fd_sc_hd__nor2_1 _0730_ (.A(net359),
    .B(_0460_),
    .Y(_0463_));
 sky130_fd_sc_hd__a31o_1 _0731_ (.A1(net359),
    .A2(_0430_),
    .A3(_0462_),
    .B1(_0463_),
    .X(_0348_));
 sky130_fd_sc_hd__a31o_1 _0732_ (.A1(net368),
    .A2(\uart_tx_inst.transmitting ),
    .A3(_0435_),
    .B1(net407),
    .X(_0464_));
 sky130_fd_sc_hd__and3_1 _0733_ (.A(_0446_),
    .B(_0460_),
    .C(net408),
    .X(_0347_));
 sky130_fd_sc_hd__or2_1 _0734_ (.A(net368),
    .B(_0435_),
    .X(_0465_));
 sky130_fd_sc_hd__a32o_1 _0735_ (.A1(_0428_),
    .A2(_0437_),
    .A3(_0465_),
    .B1(_0426_),
    .B2(net368),
    .X(_0346_));
 sky130_fd_sc_hd__a31o_1 _0736_ (.A1(\uart_tx_inst.clock_count[2] ),
    .A2(\uart_tx_inst.clock_count[1] ),
    .A3(\uart_tx_inst.clock_count[0] ),
    .B1(net315),
    .X(_0466_));
 sky130_fd_sc_hd__a32o_1 _0737_ (.A1(_0428_),
    .A2(_0436_),
    .A3(_0466_),
    .B1(_0426_),
    .B2(net315),
    .X(_0345_));
 sky130_fd_sc_hd__and3_1 _0738_ (.A(net382),
    .B(\uart_tx_inst.clock_count[0] ),
    .C(\uart_tx_inst.transmitting ),
    .X(_0467_));
 sky130_fd_sc_hd__nor2_1 _0739_ (.A(_0445_),
    .B(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__mux2_1 _0740_ (.A0(_0467_),
    .A1(_0468_),
    .S(net362),
    .X(_0344_));
 sky130_fd_sc_hd__and2_1 _0741_ (.A(\uart_tx_inst.clock_count[0] ),
    .B(\uart_tx_inst.transmitting ),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _0742_ (.A0(_0469_),
    .A1(_0468_),
    .S(net382),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _0743_ (.A0(net96),
    .A1(_0426_),
    .S(net394),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _0744_ (.A0(net220),
    .A1(net201),
    .S(\uart_tx_inst.bit_index[0] ),
    .X(_0470_));
 sky130_fd_sc_hd__nor2_1 _0745_ (.A(net388),
    .B(\uart_tx_inst.bit_index[2] ),
    .Y(_0471_));
 sky130_fd_sc_hd__a32o_1 _0746_ (.A1(net416),
    .A2(net240),
    .A3(_0471_),
    .B1(_0470_),
    .B2(net377),
    .X(_0472_));
 sky130_fd_sc_hd__and2b_1 _0747_ (.A_N(net384),
    .B(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _0748_ (.A0(net142),
    .A1(net122),
    .S(\uart_tx_inst.bit_index[0] ),
    .X(_0474_));
 sky130_fd_sc_hd__or3_1 _0749_ (.A(net377),
    .B(net384),
    .C(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__mux4_1 _0750_ (.A0(net158),
    .A1(\uart_tx_inst.shift_reg[3] ),
    .A2(net156),
    .A3(net154),
    .S0(net416),
    .S1(net377),
    .X(_0476_));
 sky130_fd_sc_hd__a22o_1 _0751_ (.A1(net388),
    .A2(_0475_),
    .B1(_0476_),
    .B2(net384),
    .X(_0477_));
 sky130_fd_sc_hd__nor2_1 _0752_ (.A(_0473_),
    .B(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__a2bb2o_1 _0753_ (.A1_N(_0478_),
    .A2_N(_0423_),
    .B1(net419),
    .B2(_0430_),
    .X(_0341_));
 sky130_fd_sc_hd__or2_1 _0754_ (.A(net122),
    .B(_0445_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _0755_ (.A0(net142),
    .A1(net130),
    .S(_0445_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _0756_ (.A0(net154),
    .A1(net120),
    .S(_0445_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _0757_ (.A0(net156),
    .A1(net140),
    .S(_0445_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _0758_ (.A0(net201),
    .A1(net128),
    .S(_0445_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _0759_ (.A0(net220),
    .A1(net124),
    .S(_0445_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _0760_ (.A0(net425),
    .A1(net134),
    .S(_0445_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _0761_ (.A0(net158),
    .A1(net136),
    .S(_0445_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _0762_ (.A0(net240),
    .A1(net138),
    .S(_0445_),
    .X(_0332_));
 sky130_fd_sc_hd__and2_2 _0763_ (.A(net97),
    .B(_0387_),
    .X(_0479_));
 sky130_fd_sc_hd__nand2_4 _0764_ (.A(net95),
    .B(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__inv_2 _0765_ (.A(_0480_),
    .Y(_0000_));
 sky130_fd_sc_hd__mux2_1 _0766_ (.A0(net181),
    .A1(net179),
    .S(_0480_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _0767_ (.A0(net144),
    .A1(\uart_rx_inst.o_data[6] ),
    .S(_0480_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _0768_ (.A0(net150),
    .A1(\uart_rx_inst.o_data[5] ),
    .S(_0480_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _0769_ (.A0(net222),
    .A1(\uart_rx_inst.o_data[4] ),
    .S(_0480_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _0770_ (.A0(net266),
    .A1(\uart_rx_inst.o_data[3] ),
    .S(_0480_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _0771_ (.A0(net183),
    .A1(\uart_rx_inst.o_data[2] ),
    .S(_0480_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _0772_ (.A0(net132),
    .A1(\uart_rx_inst.o_data[1] ),
    .S(_0480_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _0773_ (.A0(net148),
    .A1(\uart_rx_inst.o_data[0] ),
    .S(_0480_),
    .X(_0324_));
 sky130_fd_sc_hd__and2b_2 _0774_ (.A_N(net98),
    .B(net1),
    .X(_0481_));
 sky130_fd_sc_hd__nand2b_1 _0775_ (.A_N(net98),
    .B(net1),
    .Y(_0482_));
 sky130_fd_sc_hd__a21o_1 _0776_ (.A1(_0393_),
    .A2(_0482_),
    .B1(_0479_),
    .X(_0483_));
 sky130_fd_sc_hd__a221o_1 _0777_ (.A1(net97),
    .A2(net226),
    .B1(_0482_),
    .B2(_0393_),
    .C1(_0479_),
    .X(_0484_));
 sky130_fd_sc_hd__a21bo_1 _0778_ (.A1(net193),
    .A2(_0484_),
    .B1_N(_0407_),
    .X(_0323_));
 sky130_fd_sc_hd__a211oi_1 _0779_ (.A1(_0393_),
    .A2(_0482_),
    .B1(_0479_),
    .C1(_0405_),
    .Y(_0485_));
 sky130_fd_sc_hd__o21a_1 _0780_ (.A1(net225),
    .A2(_0485_),
    .B1(_0484_),
    .X(_0322_));
 sky130_fd_sc_hd__a32o_1 _0781_ (.A1(_0384_),
    .A2(_0394_),
    .A3(_0405_),
    .B1(_0483_),
    .B2(net343),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _0782_ (.A0(_0394_),
    .A1(_0483_),
    .S(net171),
    .X(_0320_));
 sky130_fd_sc_hd__nor2_1 _0783_ (.A(_0377_),
    .B(_0481_),
    .Y(_0486_));
 sky130_fd_sc_hd__and2_1 _0784_ (.A(net324),
    .B(net372),
    .X(_0487_));
 sky130_fd_sc_hd__and4_2 _0785_ (.A(net326),
    .B(net340),
    .C(net347),
    .D(net399),
    .X(_0488_));
 sky130_fd_sc_hd__nand2_1 _0786_ (.A(net380),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__and4_1 _0787_ (.A(net328),
    .B(net415),
    .C(net336),
    .D(net380),
    .X(_0490_));
 sky130_fd_sc_hd__and3_1 _0788_ (.A(net412),
    .B(_0488_),
    .C(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__and4_1 _0789_ (.A(net309),
    .B(\uart_rx_inst.clock_count[8] ),
    .C(_0488_),
    .D(_0490_),
    .X(_0492_));
 sky130_fd_sc_hd__nand2_1 _0790_ (.A(net357),
    .B(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__and3_2 _0791_ (.A(net313),
    .B(net357),
    .C(_0492_),
    .X(_0494_));
 sky130_fd_sc_hd__nand2_1 _0792_ (.A(_0487_),
    .B(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__nand3_1 _0793_ (.A(net345),
    .B(_0487_),
    .C(_0494_),
    .Y(_0496_));
 sky130_fd_sc_hd__and4_1 _0794_ (.A(net345),
    .B(net97),
    .C(_0487_),
    .D(_0494_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _0795_ (.A0(_0486_),
    .A1(_0377_),
    .S(_0497_),
    .X(_0319_));
 sky130_fd_sc_hd__nor2_2 _0796_ (.A(net1),
    .B(net98),
    .Y(_0498_));
 sky130_fd_sc_hd__a21o_1 _0797_ (.A1(_0487_),
    .A2(_0494_),
    .B1(net345),
    .X(_0499_));
 sky130_fd_sc_hd__a32o_1 _0798_ (.A1(net97),
    .A2(_0496_),
    .A3(_0499_),
    .B1(_0498_),
    .B2(net345),
    .X(_0318_));
 sky130_fd_sc_hd__nand2_1 _0799_ (.A(net372),
    .B(_0494_),
    .Y(_0500_));
 sky130_fd_sc_hd__a21o_1 _0800_ (.A1(\uart_rx_inst.clock_count[12] ),
    .A2(_0494_),
    .B1(net324),
    .X(_0501_));
 sky130_fd_sc_hd__a32o_1 _0801_ (.A1(net97),
    .A2(_0495_),
    .A3(_0501_),
    .B1(_0498_),
    .B2(net324),
    .X(_0317_));
 sky130_fd_sc_hd__or2_1 _0802_ (.A(net372),
    .B(_0494_),
    .X(_0502_));
 sky130_fd_sc_hd__and2_1 _0803_ (.A(net97),
    .B(net352),
    .X(_0503_));
 sky130_fd_sc_hd__a32o_1 _0804_ (.A1(_0500_),
    .A2(_0502_),
    .A3(_0503_),
    .B1(_0498_),
    .B2(net372),
    .X(_0316_));
 sky130_fd_sc_hd__a31o_1 _0805_ (.A1(\uart_rx_inst.clock_count[10] ),
    .A2(net98),
    .A3(_0492_),
    .B1(_0481_),
    .X(_0504_));
 sky130_fd_sc_hd__o2bb2a_1 _0806_ (.A1_N(net97),
    .A2_N(_0494_),
    .B1(_0504_),
    .B2(net313),
    .X(_0315_));
 sky130_fd_sc_hd__or2_1 _0807_ (.A(net357),
    .B(_0492_),
    .X(_0505_));
 sky130_fd_sc_hd__a32o_1 _0808_ (.A1(_0493_),
    .A2(_0503_),
    .A3(_0505_),
    .B1(_0498_),
    .B2(net357),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _0809_ (.A0(net1),
    .A1(_0491_),
    .S(net98),
    .X(_0506_));
 sky130_fd_sc_hd__o2bb2a_1 _0810_ (.A1_N(net98),
    .A2_N(_0492_),
    .B1(_0506_),
    .B2(net309),
    .X(_0313_));
 sky130_fd_sc_hd__and3_1 _0811_ (.A(_0378_),
    .B(_0488_),
    .C(_0490_),
    .X(_0507_));
 sky130_fd_sc_hd__a2bb2o_1 _0812_ (.A1_N(_0378_),
    .A2_N(_0506_),
    .B1(_0507_),
    .B2(net97),
    .X(_0312_));
 sky130_fd_sc_hd__and4_1 _0813_ (.A(net336),
    .B(net380),
    .C(net98),
    .D(_0488_),
    .X(_0508_));
 sky130_fd_sc_hd__and2_1 _0814_ (.A(net415),
    .B(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__nor2_1 _0815_ (.A(_0481_),
    .B(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__mux2_1 _0816_ (.A0(_0509_),
    .A1(_0510_),
    .S(net328),
    .X(_0311_));
 sky130_fd_sc_hd__a31o_1 _0817_ (.A1(net415),
    .A2(_0393_),
    .A3(_0482_),
    .B1(_0508_),
    .X(_0511_));
 sky130_fd_sc_hd__and2b_1 _0818_ (.A_N(_0509_),
    .B(_0511_),
    .X(_0310_));
 sky130_fd_sc_hd__a31o_1 _0819_ (.A1(\uart_rx_inst.clock_count[4] ),
    .A2(net98),
    .A3(_0488_),
    .B1(_0481_),
    .X(_0512_));
 sky130_fd_sc_hd__o21ba_1 _0820_ (.A1(net336),
    .A2(_0512_),
    .B1_N(_0508_),
    .X(_0309_));
 sky130_fd_sc_hd__or2_1 _0821_ (.A(net380),
    .B(_0488_),
    .X(_0513_));
 sky130_fd_sc_hd__a32o_1 _0822_ (.A1(_0489_),
    .A2(_0503_),
    .A3(_0513_),
    .B1(_0498_),
    .B2(net380),
    .X(_0308_));
 sky130_fd_sc_hd__and4_1 _0823_ (.A(net340),
    .B(\uart_rx_inst.clock_count[1] ),
    .C(\uart_rx_inst.clock_count[0] ),
    .D(net97),
    .X(_0514_));
 sky130_fd_sc_hd__o21ai_1 _0824_ (.A1(_0392_),
    .A2(_0488_),
    .B1(net97),
    .Y(_0515_));
 sky130_fd_sc_hd__o31a_1 _0825_ (.A1(net326),
    .A2(_0481_),
    .A3(_0514_),
    .B1(_0515_),
    .X(_0307_));
 sky130_fd_sc_hd__a31o_1 _0826_ (.A1(net347),
    .A2(\uart_rx_inst.clock_count[0] ),
    .A3(net97),
    .B1(_0481_),
    .X(_0516_));
 sky130_fd_sc_hd__o21ba_1 _0827_ (.A1(net340),
    .A2(_0516_),
    .B1_N(_0514_),
    .X(_0306_));
 sky130_fd_sc_hd__a21oi_1 _0828_ (.A1(\uart_rx_inst.clock_count[0] ),
    .A2(net97),
    .B1(net347),
    .Y(_0517_));
 sky130_fd_sc_hd__nor2_1 _0829_ (.A(_0516_),
    .B(net348),
    .Y(_0305_));
 sky130_fd_sc_hd__mux2_1 _0830_ (.A0(net97),
    .A1(_0498_),
    .S(net399),
    .X(_0304_));
 sky130_fd_sc_hd__or4b_1 _0831_ (.A(net256),
    .B(net275),
    .C(net99),
    .D_N(net210),
    .X(_0518_));
 sky130_fd_sc_hd__and2b_1 _0832_ (.A_N(net299),
    .B(net356),
    .X(_0519_));
 sky130_fd_sc_hd__and3b_2 _0833_ (.A_N(net299),
    .B(net356),
    .C(net320),
    .X(_0520_));
 sky130_fd_sc_hd__nand2_2 _0834_ (.A(net320),
    .B(_0519_),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2b_2 _0835_ (.A_N(net386),
    .B(net410),
    .Y(_0522_));
 sky130_fd_sc_hd__and3b_1 _0836_ (.A_N(_0522_),
    .B(_0518_),
    .C(_0520_),
    .X(_0523_));
 sky130_fd_sc_hd__and3b_2 _0837_ (.A_N(net418),
    .B(_0382_),
    .C(net320),
    .X(_0524_));
 sky130_fd_sc_hd__a211oi_4 _0838_ (.A1(_0520_),
    .A2(_0522_),
    .B1(_0523_),
    .C1(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__nand2b_1 _0839_ (.A_N(net422),
    .B(net99),
    .Y(_0526_));
 sky130_fd_sc_hd__or2_4 _0840_ (.A(net210),
    .B(net275),
    .X(_0527_));
 sky130_fd_sc_hd__or4b_2 _0841_ (.A(net256),
    .B(net210),
    .C(net342),
    .D_N(net99),
    .X(_0528_));
 sky130_fd_sc_hd__and2b_1 _0842_ (.A_N(net320),
    .B(_0519_),
    .X(_0529_));
 sky130_fd_sc_hd__and4bb_4 _0843_ (.A_N(net421),
    .B_N(net423),
    .C(net247),
    .D(net418),
    .X(_0530_));
 sky130_fd_sc_hd__and2b_1 _0844_ (.A_N(net320),
    .B(net356),
    .X(_0531_));
 sky130_fd_sc_hd__and3b_2 _0845_ (.A_N(net320),
    .B(net356),
    .C(net299),
    .X(_0532_));
 sky130_fd_sc_hd__o31a_1 _0846_ (.A1(net210),
    .A2(_0381_),
    .A3(_0526_),
    .B1(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__and2b_1 _0847_ (.A_N(net247),
    .B(_0531_),
    .X(_0534_));
 sky130_fd_sc_hd__a211oi_2 _0848_ (.A1(_0528_),
    .A2(_0530_),
    .B1(_0533_),
    .C1(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__nor3_1 _0849_ (.A(net421),
    .B(net418),
    .C(net299),
    .Y(_0536_));
 sky130_fd_sc_hd__or3_2 _0850_ (.A(net320),
    .B(net356),
    .C(net299),
    .X(_0537_));
 sky130_fd_sc_hd__o211a_1 _0851_ (.A1(net247),
    .A2(_0537_),
    .B1(_0535_),
    .C1(_0525_),
    .X(_0538_));
 sky130_fd_sc_hd__and3b_1 _0852_ (.A_N(net356),
    .B(net299),
    .C(net320),
    .X(_0539_));
 sky130_fd_sc_hd__and4b_1 _0853_ (.A_N(net301),
    .B(net306),
    .C(net285),
    .D(net305),
    .X(_0540_));
 sky130_fd_sc_hd__and4b_1 _0854_ (.A_N(net311),
    .B(net304),
    .C(net323),
    .D(net292),
    .X(_0541_));
 sky130_fd_sc_hd__nand2_1 _0855_ (.A(_0540_),
    .B(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__and3_1 _0856_ (.A(_0529_),
    .B(_0540_),
    .C(_0541_),
    .X(_0543_));
 sky130_fd_sc_hd__or3_1 _0857_ (.A(net321),
    .B(_0539_),
    .C(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__a21bo_1 _0858_ (.A1(_0538_),
    .A2(_0544_),
    .B1_N(_0525_),
    .X(_0303_));
 sky130_fd_sc_hd__and4bb_1 _0859_ (.A_N(net304),
    .B_N(net292),
    .C(net323),
    .D(net311),
    .X(_0545_));
 sky130_fd_sc_hd__and4bb_1 _0860_ (.A_N(net306),
    .B_N(net305),
    .C(net285),
    .D(net301),
    .X(_0546_));
 sky130_fd_sc_hd__a31o_1 _0861_ (.A1(_0529_),
    .A2(_0545_),
    .A3(_0546_),
    .B1(_0539_),
    .X(_0547_));
 sky130_fd_sc_hd__or4b_1 _0862_ (.A(\uart_rx_inst.o_data[4] ),
    .B(\uart_rx_inst.o_data[2] ),
    .C(\uart_rx_inst.o_data[0] ),
    .D_N(\uart_rx_inst.o_data[3] ),
    .X(_0548_));
 sky130_fd_sc_hd__nor3_1 _0863_ (.A(_0373_),
    .B(net281),
    .C(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__and4b_1 _0864_ (.A_N(\uart_rx_inst.o_data[3] ),
    .B(net286),
    .C(net228),
    .D(net288),
    .X(_0550_));
 sky130_fd_sc_hd__a31o_1 _0865_ (.A1(_0373_),
    .A2(net281),
    .A3(_0550_),
    .B1(_0549_),
    .X(_0551_));
 sky130_fd_sc_hd__a41o_1 _0866_ (.A1(net263),
    .A2(net169),
    .A3(net300),
    .A4(_0551_),
    .B1(_0547_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _0867_ (.A0(net356),
    .A1(_0552_),
    .S(_0538_),
    .X(_0302_));
 sky130_fd_sc_hd__a21oi_1 _0868_ (.A1(_0525_),
    .A2(_0535_),
    .B1(_0379_),
    .Y(_0553_));
 sky130_fd_sc_hd__a21bo_1 _0869_ (.A1(_0545_),
    .A2(_0546_),
    .B1_N(_0542_),
    .X(_0554_));
 sky130_fd_sc_hd__a31o_1 _0870_ (.A1(_0529_),
    .A2(_0538_),
    .A3(_0554_),
    .B1(_0553_),
    .X(_0301_));
 sky130_fd_sc_hd__nor4_1 _0871_ (.A(_0519_),
    .B(_0532_),
    .C(_0536_),
    .D(_0539_),
    .Y(_0555_));
 sky130_fd_sc_hd__a2bb2o_2 _0872_ (.A1_N(net247),
    .A2_N(_0537_),
    .B1(_0522_),
    .B2(_0520_),
    .X(_0556_));
 sky130_fd_sc_hd__a2111oi_4 _0873_ (.A1(net299),
    .A2(_0524_),
    .B1(_0534_),
    .C1(net94),
    .D1(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__nor2_1 _0874_ (.A(_0520_),
    .B(_0532_),
    .Y(_0558_));
 sky130_fd_sc_hd__and3b_1 _0875_ (.A_N(_0529_),
    .B(_0557_),
    .C(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__and2_1 _0876_ (.A(net275),
    .B(net99),
    .X(_0560_));
 sky130_fd_sc_hd__nand3_1 _0877_ (.A(net210),
    .B(_0557_),
    .C(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__a31o_1 _0878_ (.A1(net210),
    .A2(_0557_),
    .A3(_0560_),
    .B1(_0380_),
    .X(_0562_));
 sky130_fd_sc_hd__nand4_1 _0879_ (.A(_0380_),
    .B(net210),
    .C(_0557_),
    .D(_0560_),
    .Y(_0563_));
 sky130_fd_sc_hd__a21oi_1 _0880_ (.A1(_0562_),
    .A2(_0563_),
    .B1(_0559_),
    .Y(_0300_));
 sky130_fd_sc_hd__a21o_1 _0881_ (.A1(_0557_),
    .A2(_0560_),
    .B1(net210),
    .X(_0564_));
 sky130_fd_sc_hd__and3b_1 _0882_ (.A_N(_0559_),
    .B(_0561_),
    .C(_0564_),
    .X(_0299_));
 sky130_fd_sc_hd__and2_1 _0883_ (.A(net99),
    .B(_0557_),
    .X(_0565_));
 sky130_fd_sc_hd__nand2_1 _0884_ (.A(_0528_),
    .B(_0529_),
    .Y(_0566_));
 sky130_fd_sc_hd__a21o_1 _0885_ (.A1(_0558_),
    .A2(_0566_),
    .B1(_0560_),
    .X(_0567_));
 sky130_fd_sc_hd__o2bb2a_1 _0886_ (.A1_N(_0557_),
    .A2_N(_0567_),
    .B1(_0565_),
    .B2(net275),
    .X(_0298_));
 sky130_fd_sc_hd__a21o_1 _0887_ (.A1(net356),
    .A2(_0557_),
    .B1(net99),
    .X(_0568_));
 sky130_fd_sc_hd__and2b_1 _0888_ (.A_N(_0565_),
    .B(_0568_),
    .X(_0297_));
 sky130_fd_sc_hd__and2_4 _0889_ (.A(net247),
    .B(_0532_),
    .X(_0569_));
 sky130_fd_sc_hd__or3b_4 _0890_ (.A(net210),
    .B(_0381_),
    .C_N(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__or3_1 _0891_ (.A(_0373_),
    .B(\byte_count[3] ),
    .C(net205),
    .X(_0571_));
 sky130_fd_sc_hd__nand2_1 _0892_ (.A(net247),
    .B(_0536_),
    .Y(_0572_));
 sky130_fd_sc_hd__a2bb2o_1 _0893_ (.A1_N(_0570_),
    .A2_N(net206),
    .B1(net92),
    .B2(net199),
    .X(_0296_));
 sky130_fd_sc_hd__or3b_1 _0894_ (.A(net256),
    .B(net205),
    .C_N(net281),
    .X(_0573_));
 sky130_fd_sc_hd__a2bb2o_1 _0895_ (.A1_N(_0570_),
    .A2_N(_0573_),
    .B1(net91),
    .B2(net273),
    .X(_0295_));
 sky130_fd_sc_hd__or3b_1 _0896_ (.A(net256),
    .B(net99),
    .C_N(net263),
    .X(_0574_));
 sky130_fd_sc_hd__a2bb2o_1 _0897_ (.A1_N(_0570_),
    .A2_N(_0574_),
    .B1(net93),
    .B2(net294),
    .X(_0294_));
 sky130_fd_sc_hd__or3b_1 _0898_ (.A(net256),
    .B(net99),
    .C_N(net288),
    .X(_0575_));
 sky130_fd_sc_hd__a2bb2o_1 _0899_ (.A1_N(_0570_),
    .A2_N(_0575_),
    .B1(net93),
    .B2(net118),
    .X(_0293_));
 sky130_fd_sc_hd__or3b_1 _0900_ (.A(net256),
    .B(net99),
    .C_N(net277),
    .X(_0576_));
 sky130_fd_sc_hd__a2bb2o_1 _0901_ (.A1_N(_0570_),
    .A2_N(_0576_),
    .B1(net92),
    .B2(net271),
    .X(_0292_));
 sky130_fd_sc_hd__or3b_1 _0902_ (.A(net256),
    .B(net99),
    .C_N(\uart_rx_inst.o_data[2] ),
    .X(_0577_));
 sky130_fd_sc_hd__a2bb2o_1 _0903_ (.A1_N(_0570_),
    .A2_N(net257),
    .B1(net92),
    .B2(net250),
    .X(_0291_));
 sky130_fd_sc_hd__or3b_1 _0904_ (.A(net256),
    .B(net205),
    .C_N(net169),
    .X(_0578_));
 sky130_fd_sc_hd__a2bb2o_1 _0905_ (.A1_N(_0570_),
    .A2_N(_0578_),
    .B1(net92),
    .B2(net254),
    .X(_0290_));
 sky130_fd_sc_hd__or3b_1 _0906_ (.A(net256),
    .B(net205),
    .C_N(net228),
    .X(_0579_));
 sky130_fd_sc_hd__a2bb2o_1 _0907_ (.A1_N(_0570_),
    .A2_N(_0579_),
    .B1(net93),
    .B2(net126),
    .X(_0289_));
 sky130_fd_sc_hd__and2b_4 _0908_ (.A_N(_0528_),
    .B(_0569_),
    .X(_0580_));
 sky130_fd_sc_hd__a22o_1 _0909_ (.A1(net218),
    .A2(net93),
    .B1(_0580_),
    .B2(net179),
    .X(_0288_));
 sky130_fd_sc_hd__a22o_1 _0910_ (.A1(net177),
    .A2(net93),
    .B1(_0580_),
    .B2(\uart_rx_inst.o_data[6] ),
    .X(_0287_));
 sky130_fd_sc_hd__a22o_1 _0911_ (.A1(net290),
    .A2(net91),
    .B1(_0580_),
    .B2(net263),
    .X(_0286_));
 sky130_fd_sc_hd__a22o_1 _0912_ (.A1(net242),
    .A2(net91),
    .B1(_0580_),
    .B2(\uart_rx_inst.o_data[4] ),
    .X(_0285_));
 sky130_fd_sc_hd__a22o_1 _0913_ (.A1(net152),
    .A2(net93),
    .B1(_0580_),
    .B2(\uart_rx_inst.o_data[3] ),
    .X(_0284_));
 sky130_fd_sc_hd__a22o_1 _0914_ (.A1(net185),
    .A2(net93),
    .B1(_0580_),
    .B2(net286),
    .X(_0283_));
 sky130_fd_sc_hd__a22o_1 _0915_ (.A1(net116),
    .A2(net93),
    .B1(_0580_),
    .B2(net169),
    .X(_0282_));
 sky130_fd_sc_hd__a22o_1 _0916_ (.A1(net252),
    .A2(net93),
    .B1(_0580_),
    .B2(net228),
    .X(_0281_));
 sky130_fd_sc_hd__nor2_1 _0917_ (.A(_0527_),
    .B(net206),
    .Y(_0581_));
 sky130_fd_sc_hd__a22o_1 _0918_ (.A1(net261),
    .A2(net92),
    .B1(_0581_),
    .B2(_0569_),
    .X(_0280_));
 sky130_fd_sc_hd__nor2_1 _0919_ (.A(_0527_),
    .B(_0573_),
    .Y(_0582_));
 sky130_fd_sc_hd__a22o_1 _0920_ (.A1(net297),
    .A2(net91),
    .B1(_0582_),
    .B2(_0569_),
    .X(_0279_));
 sky130_fd_sc_hd__nor2_1 _0921_ (.A(_0527_),
    .B(_0574_),
    .Y(_0583_));
 sky130_fd_sc_hd__a22o_1 _0922_ (.A1(net160),
    .A2(net92),
    .B1(net264),
    .B2(_0569_),
    .X(_0278_));
 sky130_fd_sc_hd__nor2_1 _0923_ (.A(_0527_),
    .B(_0575_),
    .Y(_0584_));
 sky130_fd_sc_hd__a22o_1 _0924_ (.A1(net307),
    .A2(net92),
    .B1(_0584_),
    .B2(_0569_),
    .X(_0277_));
 sky130_fd_sc_hd__nor2_1 _0925_ (.A(_0527_),
    .B(_0576_),
    .Y(_0585_));
 sky130_fd_sc_hd__a22o_1 _0926_ (.A1(net338),
    .A2(net92),
    .B1(_0585_),
    .B2(_0569_),
    .X(_0276_));
 sky130_fd_sc_hd__nor2_1 _0927_ (.A(_0527_),
    .B(net257),
    .Y(_0586_));
 sky130_fd_sc_hd__a22o_1 _0928_ (.A1(net375),
    .A2(net91),
    .B1(_0586_),
    .B2(_0569_),
    .X(_0275_));
 sky130_fd_sc_hd__nor2_1 _0929_ (.A(_0527_),
    .B(_0578_),
    .Y(_0587_));
 sky130_fd_sc_hd__a22o_1 _0930_ (.A1(net317),
    .A2(net91),
    .B1(_0587_),
    .B2(net322),
    .X(_0274_));
 sky130_fd_sc_hd__nor2_1 _0931_ (.A(_0527_),
    .B(_0579_),
    .Y(_0588_));
 sky130_fd_sc_hd__a22o_1 _0932_ (.A1(net233),
    .A2(net91),
    .B1(_0588_),
    .B2(_0569_),
    .X(_0273_));
 sky130_fd_sc_hd__and2b_4 _0933_ (.A_N(_0528_),
    .B(_0530_),
    .X(_0589_));
 sky130_fd_sc_hd__a22o_1 _0934_ (.A1(net175),
    .A2(net93),
    .B1(_0589_),
    .B2(net179),
    .X(_0272_));
 sky130_fd_sc_hd__a22o_1 _0935_ (.A1(net259),
    .A2(net92),
    .B1(_0589_),
    .B2(\uart_rx_inst.o_data[6] ),
    .X(_0271_));
 sky130_fd_sc_hd__a22o_1 _0936_ (.A1(net187),
    .A2(net93),
    .B1(_0589_),
    .B2(\uart_rx_inst.o_data[5] ),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_1 _0937_ (.A1(net229),
    .A2(net91),
    .B1(_0589_),
    .B2(\uart_rx_inst.o_data[4] ),
    .X(_0269_));
 sky130_fd_sc_hd__a22o_1 _0938_ (.A1(net165),
    .A2(net93),
    .B1(_0589_),
    .B2(\uart_rx_inst.o_data[3] ),
    .X(_0268_));
 sky130_fd_sc_hd__a22o_1 _0939_ (.A1(net231),
    .A2(net92),
    .B1(_0589_),
    .B2(\uart_rx_inst.o_data[2] ),
    .X(_0267_));
 sky130_fd_sc_hd__a22o_1 _0940_ (.A1(net167),
    .A2(net93),
    .B1(_0589_),
    .B2(\uart_rx_inst.o_data[1] ),
    .X(_0266_));
 sky130_fd_sc_hd__a22o_1 _0941_ (.A1(net146),
    .A2(net92),
    .B1(_0589_),
    .B2(net228),
    .X(_0265_));
 sky130_fd_sc_hd__a22o_1 _0942_ (.A1(net280),
    .A2(net91),
    .B1(_0581_),
    .B2(net248),
    .X(_0264_));
 sky130_fd_sc_hd__a22o_1 _0943_ (.A1(net269),
    .A2(net92),
    .B1(_0582_),
    .B2(net248),
    .X(_0263_));
 sky130_fd_sc_hd__a22o_1 _0944_ (.A1(net191),
    .A2(net92),
    .B1(_0583_),
    .B2(net248),
    .X(_0262_));
 sky130_fd_sc_hd__a22o_1 _0945_ (.A1(net189),
    .A2(net93),
    .B1(_0584_),
    .B2(_0530_),
    .X(_0261_));
 sky130_fd_sc_hd__a22o_1 _0946_ (.A1(net216),
    .A2(net93),
    .B1(_0585_),
    .B2(_0530_),
    .X(_0260_));
 sky130_fd_sc_hd__a22o_1 _0947_ (.A1(net244),
    .A2(net92),
    .B1(_0586_),
    .B2(_0530_),
    .X(_0259_));
 sky130_fd_sc_hd__a22o_1 _0948_ (.A1(net330),
    .A2(net92),
    .B1(_0587_),
    .B2(net248),
    .X(_0258_));
 sky130_fd_sc_hd__a22o_1 _0949_ (.A1(net208),
    .A2(_0572_),
    .B1(_0588_),
    .B2(_0530_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _0950_ (.A0(net179),
    .A1(net301),
    .S(net91),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _0951_ (.A0(net281),
    .A1(net306),
    .S(net91),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _0952_ (.A0(net263),
    .A1(net285),
    .S(net91),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _0953_ (.A0(net288),
    .A1(net305),
    .S(net91),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _0954_ (.A0(net277),
    .A1(net311),
    .S(net91),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _0955_ (.A0(net286),
    .A1(net304),
    .S(net91),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _0956_ (.A0(net169),
    .A1(net323),
    .S(net91),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _0957_ (.A0(net228),
    .A1(net292),
    .S(_0572_),
    .X(_0249_));
 sky130_fd_sc_hd__a21o_4 _0958_ (.A1(_0521_),
    .A2(_0537_),
    .B1(_0556_),
    .X(_0590_));
 sky130_fd_sc_hd__nor3_4 _0959_ (.A(\byte_count[3] ),
    .B(net210),
    .C(_0521_),
    .Y(_0591_));
 sky130_fd_sc_hd__mux4_1 _0960_ (.A0(net34),
    .A1(net11),
    .A2(net20),
    .A3(net29),
    .S0(net99),
    .S1(\byte_count[1] ),
    .X(_0592_));
 sky130_fd_sc_hd__and3b_1 _0961_ (.A_N(_0590_),
    .B(_0591_),
    .C(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__a21o_1 _0962_ (.A1(net130),
    .A2(_0590_),
    .B1(_0593_),
    .X(_0248_));
 sky130_fd_sc_hd__mux4_1 _0963_ (.A0(net33),
    .A1(net10),
    .A2(net19),
    .A3(net28),
    .S0(net99),
    .S1(\byte_count[1] ),
    .X(_0594_));
 sky130_fd_sc_hd__and3b_1 _0964_ (.A_N(_0590_),
    .B(_0591_),
    .C(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__a21o_1 _0965_ (.A1(net120),
    .A2(_0590_),
    .B1(_0595_),
    .X(_0247_));
 sky130_fd_sc_hd__mux4_1 _0966_ (.A0(net32),
    .A1(net9),
    .A2(net18),
    .A3(net26),
    .S0(net99),
    .S1(\byte_count[1] ),
    .X(_0596_));
 sky130_fd_sc_hd__and3b_1 _0967_ (.A_N(_0590_),
    .B(_0591_),
    .C(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__a21o_1 _0968_ (.A1(net140),
    .A2(_0590_),
    .B1(_0597_),
    .X(_0246_));
 sky130_fd_sc_hd__mux4_1 _0969_ (.A0(net31),
    .A1(net8),
    .A2(net17),
    .A3(net25),
    .S0(\byte_count[0] ),
    .S1(\byte_count[1] ),
    .X(_0598_));
 sky130_fd_sc_hd__and3b_1 _0970_ (.A_N(_0590_),
    .B(_0591_),
    .C(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__a21o_1 _0971_ (.A1(net128),
    .A2(_0590_),
    .B1(_0599_),
    .X(_0245_));
 sky130_fd_sc_hd__mux4_1 _0972_ (.A0(net30),
    .A1(net7),
    .A2(net15),
    .A3(net24),
    .S0(net99),
    .S1(\byte_count[1] ),
    .X(_0600_));
 sky130_fd_sc_hd__and3b_1 _0973_ (.A_N(_0590_),
    .B(_0591_),
    .C(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__a21o_1 _0974_ (.A1(net124),
    .A2(_0590_),
    .B1(_0601_),
    .X(_0244_));
 sky130_fd_sc_hd__mux4_1 _0975_ (.A0(net27),
    .A1(net6),
    .A2(net14),
    .A3(net23),
    .S0(net99),
    .S1(\byte_count[1] ),
    .X(_0602_));
 sky130_fd_sc_hd__and3b_1 _0976_ (.A_N(_0590_),
    .B(net211),
    .C(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__a21o_1 _0977_ (.A1(net134),
    .A2(_0590_),
    .B1(net212),
    .X(_0243_));
 sky130_fd_sc_hd__mux4_1 _0978_ (.A0(net16),
    .A1(net36),
    .A2(net13),
    .A3(net22),
    .S0(net99),
    .S1(\byte_count[1] ),
    .X(_0604_));
 sky130_fd_sc_hd__and3b_1 _0979_ (.A_N(_0590_),
    .B(_0591_),
    .C(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__a21o_1 _0980_ (.A1(net136),
    .A2(_0590_),
    .B1(_0605_),
    .X(_0242_));
 sky130_fd_sc_hd__mux4_1 _0981_ (.A0(net5),
    .A1(net35),
    .A2(net12),
    .A3(net21),
    .S0(\byte_count[0] ),
    .S1(\byte_count[1] ),
    .X(_0606_));
 sky130_fd_sc_hd__and3b_1 _0982_ (.A_N(_0590_),
    .B(_0591_),
    .C(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__a21o_1 _0983_ (.A1(net138),
    .A2(_0590_),
    .B1(_0607_),
    .X(_0241_));
 sky130_fd_sc_hd__a31o_1 _0984_ (.A1(net386),
    .A2(_0521_),
    .A3(_0537_),
    .B1(_0523_),
    .X(_0240_));
 sky130_fd_sc_hd__nand2_1 _0985_ (.A(_0542_),
    .B(_0589_),
    .Y(_0608_));
 sky130_fd_sc_hd__o21ai_1 _0986_ (.A1(net356),
    .A2(_0382_),
    .B1(net320),
    .Y(_0609_));
 sky130_fd_sc_hd__a211o_1 _0987_ (.A1(net356),
    .A2(net247),
    .B1(_0379_),
    .C1(net320),
    .X(_0610_));
 sky130_fd_sc_hd__and4_1 _0988_ (.A(_0535_),
    .B(_0608_),
    .C(_0609_),
    .D(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__nor2_2 _0989_ (.A(_0526_),
    .B(_0570_),
    .Y(_0612_));
 sky130_fd_sc_hd__mux2_1 _0990_ (.A0(net361),
    .A1(net179),
    .S(net89),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _0991_ (.A0(net370),
    .A1(net281),
    .S(net90),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _0992_ (.A0(net374),
    .A1(net263),
    .S(net90),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _0993_ (.A0(net365),
    .A1(net288),
    .S(net89),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _0994_ (.A0(net390),
    .A1(net277),
    .S(net89),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _0995_ (.A0(net373),
    .A1(net286),
    .S(net90),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(net364),
    .A1(net169),
    .S(net89),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _0997_ (.A0(net379),
    .A1(net228),
    .S(net90),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _0998_ (.A0(net70),
    .A1(net199),
    .S(net89),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _0999_ (.A0(net69),
    .A1(net273),
    .S(net89),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _1000_ (.A0(net68),
    .A1(net294),
    .S(net90),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _1001_ (.A0(net67),
    .A1(net118),
    .S(net90),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _1002_ (.A0(net65),
    .A1(net271),
    .S(net89),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _1003_ (.A0(net64),
    .A1(net250),
    .S(_0612_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _1004_ (.A0(net63),
    .A1(net254),
    .S(net89),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _1005_ (.A0(net62),
    .A1(net126),
    .S(net90),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _1006_ (.A0(net246),
    .A1(net218),
    .S(net90),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _1007_ (.A0(net224),
    .A1(net177),
    .S(net90),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _1008_ (.A0(net59),
    .A1(net290),
    .S(net89),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _1009_ (.A0(net279),
    .A1(net242),
    .S(net89),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _1010_ (.A0(net195),
    .A1(net152),
    .S(net90),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _1011_ (.A0(net56),
    .A1(net185),
    .S(net90),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _1012_ (.A0(net86),
    .A1(net116),
    .S(net90),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _1013_ (.A0(net283),
    .A1(net252),
    .S(net90),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _1014_ (.A0(net284),
    .A1(net261),
    .S(net89),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _1015_ (.A0(net312),
    .A1(net297),
    .S(net89),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _1016_ (.A0(net82),
    .A1(net160),
    .S(net89),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _1017_ (.A0(net319),
    .A1(net307),
    .S(net89),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _1018_ (.A0(net80),
    .A1(net338),
    .S(net90),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _1019_ (.A0(net77),
    .A1(net375),
    .S(net90),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _1020_ (.A0(net66),
    .A1(net317),
    .S(net89),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _1021_ (.A0(net276),
    .A1(net233),
    .S(net89),
    .X(_0208_));
 sky130_fd_sc_hd__o2bb2a_1 _1022_ (.A1_N(_0528_),
    .A2_N(_0530_),
    .B1(_0531_),
    .B2(_0379_),
    .X(_0613_));
 sky130_fd_sc_hd__a21boi_1 _1023_ (.A1(_0542_),
    .A2(_0589_),
    .B1_N(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__and3_1 _1024_ (.A(_0525_),
    .B(_0535_),
    .C(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__and4_4 _1025_ (.A(_0525_),
    .B(_0531_),
    .C(_0535_),
    .D(_0614_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _1026_ (.A0(net44),
    .A1(net175),
    .S(_0616_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _1027_ (.A0(net278),
    .A1(net259),
    .S(_0616_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _1028_ (.A0(net214),
    .A1(net187),
    .S(_0616_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _1029_ (.A0(net238),
    .A1(net229),
    .S(_0616_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _1030_ (.A0(net197),
    .A1(net165),
    .S(_0616_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _1031_ (.A0(net265),
    .A1(net231),
    .S(_0616_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _1032_ (.A0(net203),
    .A1(net167),
    .S(_0616_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _1033_ (.A0(net52),
    .A1(net146),
    .S(_0616_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _1034_ (.A0(net296),
    .A1(net280),
    .S(_0616_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _1035_ (.A0(net289),
    .A1(net269),
    .S(_0616_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _1036_ (.A0(net49),
    .A1(net191),
    .S(_0616_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _1037_ (.A0(net235),
    .A1(net189),
    .S(_0616_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _1038_ (.A0(net282),
    .A1(net216),
    .S(_0616_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _1039_ (.A0(net268),
    .A1(net244),
    .S(_0616_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _1040_ (.A0(net335),
    .A1(net330),
    .S(_0616_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _1041_ (.A0(net236),
    .A1(net208),
    .S(_0616_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _1042_ (.A0(net371),
    .A1(net321),
    .S(_0611_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _1043_ (.A0(net417),
    .A1(_0531_),
    .S(_0615_),
    .X(_0190_));
 sky130_fd_sc_hd__o2111a_1 _1044_ (.A1(net377),
    .A2(net384),
    .B1(net96),
    .C1(_0422_),
    .D1(net388),
    .X(_0370_));
 sky130_fd_sc_hd__a21o_1 _1045_ (.A1(net410),
    .A2(_0446_),
    .B1(_0370_),
    .X(_0189_));
 sky130_fd_sc_hd__and2b_1 _1046_ (.A_N(net162),
    .B(net1),
    .X(_0371_));
 sky130_fd_sc_hd__o21a_1 _1047_ (.A1(net98),
    .A2(_0371_),
    .B1(_0480_),
    .X(_0001_));
 sky130_fd_sc_hd__nor2_1 _1048_ (.A(_0426_),
    .B(_0370_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _1049_ (.A(net111),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _1050_ (.A(net104),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _1051_ (.A(net109),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _1052_ (.A(net112),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _1053_ (.A(net109),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _1054_ (.A(net111),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _1055_ (.A(net101),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _1056_ (.A(net112),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _1057_ (.A(net109),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _1058_ (.A(net107),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1059_ (.A(net112),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _1060_ (.A(net104),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _1061_ (.A(net109),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(net104),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _1063_ (.A(net107),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _1064_ (.A(net101),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _1065_ (.A(net109),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _1066_ (.A(net100),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _1067_ (.A(net107),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _1068_ (.A(net107),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _1069_ (.A(net100),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1070_ (.A(net100),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _1071_ (.A(net109),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1072_ (.A(net112),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1073_ (.A(net109),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1074_ (.A(net109),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _1075_ (.A(net102),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _1076_ (.A(net101),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _1077_ (.A(net103),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _1078_ (.A(net101),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1079_ (.A(net107),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _1080_ (.A(net109),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1081_ (.A(net100),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _1082_ (.A(net100),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _1083_ (.A(net100),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _1084_ (.A(net110),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1085_ (.A(net112),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _1086_ (.A(net112),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _1087_ (.A(net101),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _1088_ (.A(net100),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _1089_ (.A(net110),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _1090_ (.A(net110),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _1091_ (.A(net100),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _1092_ (.A(net112),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _1093_ (.A(net103),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _1094_ (.A(net109),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _1095_ (.A(net104),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _1096_ (.A(net100),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _1097_ (.A(net101),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _1098_ (.A(net111),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _1099_ (.A(net101),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _1100_ (.A(net104),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _1101_ (.A(net102),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _1102_ (.A(net100),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _1103_ (.A(net100),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _1104_ (.A(net104),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _1105_ (.A(net100),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _1106_ (.A(net100),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _1107_ (.A(net102),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _1108_ (.A(net108),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _1109_ (.A(net107),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _1110_ (.A(net108),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _1111_ (.A(net107),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _1112_ (.A(net107),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _1113_ (.A(net107),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _1114_ (.A(net107),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _1115_ (.A(net107),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _1116_ (.A(net110),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _1117_ (.A(net110),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _1118_ (.A(net109),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _1119_ (.A(net108),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _1120_ (.A(net101),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _1121_ (.A(net112),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _1122_ (.A(net109),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _1123_ (.A(net107),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _1124_ (.A(net112),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _1125_ (.A(net104),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _1126_ (.A(net110),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _1127_ (.A(net104),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _1128_ (.A(net107),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _1129_ (.A(net101),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _1130_ (.A(net109),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _1131_ (.A(net101),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _1132_ (.A(net107),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _1133_ (.A(net109),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _1134_ (.A(net108),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _1135_ (.A(net108),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _1136_ (.A(net110),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _1137_ (.A(net112),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _1138_ (.A(net109),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _1139_ (.A(net109),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _1140_ (.A(net102),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _1141_ (.A(net101),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _1142_ (.A(net102),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _1143_ (.A(net101),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _1144_ (.A(net107),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _1145_ (.A(net107),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _1146_ (.A(net100),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _1147_ (.A(net100),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _1148_ (.A(net106),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _1149_ (.A(net110),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _1150_ (.A(net110),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _1151_ (.A(net110),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _1152_ (.A(net101),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _1153_ (.A(net100),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _1154_ (.A(net110),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _1155_ (.A(net110),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _1156_ (.A(net101),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _1157_ (.A(net101),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _1158_ (.A(net101),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _1159_ (.A(net106),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _1160_ (.A(net108),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _1161_ (.A(net108),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _1162_ (.A(net108),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _1163_ (.A(net104),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _1164_ (.A(net111),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _1165_ (.A(net112),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _1166_ (.A(net112),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _1167_ (.A(net112),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _1168_ (.A(net112),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _1169_ (.A(net113),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _1170_ (.A(net113),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _1171_ (.A(net113),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _1172_ (.A(net113),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _1173_ (.A(net113),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _1174_ (.A(net113),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _1175_ (.A(net113),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _1176_ (.A(net113),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _1177_ (.A(net113),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _1178_ (.A(net113),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _1179_ (.A(net112),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _1180_ (.A(net112),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _1181_ (.A(net111),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _1182_ (.A(net114),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _1183_ (.A(net114),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _1184_ (.A(net111),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _1185_ (.A(net111),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _1186_ (.A(net111),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _1187_ (.A(net114),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _1188_ (.A(net111),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _1189_ (.A(net114),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _1190_ (.A(net111),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _1191_ (.A(net111),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _1192_ (.A(net104),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _1193_ (.A(net111),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _1194_ (.A(net104),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _1195_ (.A(net102),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _1196_ (.A(net102),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _1197_ (.A(net106),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _1198_ (.A(net104),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _1199_ (.A(net102),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _1200_ (.A(net102),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _1201_ (.A(net102),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _1202_ (.A(net102),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _1203_ (.A(net104),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _1204_ (.A(net104),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _1205_ (.A(net102),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _1206_ (.A(net105),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _1207_ (.A(net105),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _1208_ (.A(net105),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _1209_ (.A(net105),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _1210_ (.A(net105),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _1211_ (.A(net105),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _1212_ (.A(net103),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _1213_ (.A(net103),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _1214_ (.A(net103),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _1215_ (.A(net103),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _1216_ (.A(net103),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _1217_ (.A(net103),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _1218_ (.A(net103),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _1219_ (.A(net105),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _1220_ (.A(net105),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _1221_ (.A(net105),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _1222_ (.A(net102),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _1223_ (.A(net102),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _1224_ (.A(net102),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _1225_ (.A(net102),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _1226_ (.A(net111),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _1227_ (.A(net111),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _1228_ (.A(net114),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _1229_ (.A(net111),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _1230_ (.A(net114),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _1231_ (.A(net104),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _1232_ (.A(net111),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _1233_ (.A(net114),
    .Y(_0188_));
 sky130_fd_sc_hd__dfstp_1 _1234_ (.CLK(clknet_4_9_0_clk),
    .D(net411),
    .SET_B(_0003_),
    .Q(\uart_tx_inst.o_ready ));
 sky130_fd_sc_hd__dfrtp_4 _1235_ (.CLK(clknet_4_6_0_clk),
    .D(_0190_),
    .RESET_B(_0004_),
    .Q(net54));
 sky130_fd_sc_hd__dfrtp_2 _1236_ (.CLK(clknet_4_9_0_clk),
    .D(_0191_),
    .RESET_B(_0005_),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_1 _1237_ (.CLK(clknet_4_6_0_clk),
    .D(net237),
    .RESET_B(_0006_),
    .Q(net38));
 sky130_fd_sc_hd__dfrtp_2 _1238_ (.CLK(clknet_4_13_0_clk),
    .D(_0193_),
    .RESET_B(_0007_),
    .Q(net45));
 sky130_fd_sc_hd__dfrtp_1 _1239_ (.CLK(clknet_4_5_0_clk),
    .D(_0194_),
    .RESET_B(_0008_),
    .Q(net46));
 sky130_fd_sc_hd__dfrtp_2 _1240_ (.CLK(clknet_4_6_0_clk),
    .D(_0195_),
    .RESET_B(_0009_),
    .Q(net47));
 sky130_fd_sc_hd__dfrtp_2 _1241_ (.CLK(clknet_4_1_0_clk),
    .D(_0196_),
    .RESET_B(_0010_),
    .Q(net48));
 sky130_fd_sc_hd__dfrtp_2 _1242_ (.CLK(clknet_4_13_0_clk),
    .D(net192),
    .RESET_B(_0011_),
    .Q(net49));
 sky130_fd_sc_hd__dfrtp_1 _1243_ (.CLK(clknet_4_5_0_clk),
    .D(_0198_),
    .RESET_B(_0012_),
    .Q(net50));
 sky130_fd_sc_hd__dfrtp_1 _1244_ (.CLK(clknet_4_4_0_clk),
    .D(_0199_),
    .RESET_B(_0013_),
    .Q(net51));
 sky130_fd_sc_hd__dfrtp_2 _1245_ (.CLK(clknet_4_13_0_clk),
    .D(net147),
    .RESET_B(_0014_),
    .Q(net52));
 sky130_fd_sc_hd__dfrtp_2 _1246_ (.CLK(clknet_4_9_0_clk),
    .D(net204),
    .RESET_B(_0015_),
    .Q(net53));
 sky130_fd_sc_hd__dfrtp_1 _1247_ (.CLK(clknet_4_7_0_clk),
    .D(_0202_),
    .RESET_B(_0016_),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_2 _1248_ (.CLK(clknet_4_9_0_clk),
    .D(net198),
    .RESET_B(_0017_),
    .Q(net40));
 sky130_fd_sc_hd__dfrtp_2 _1249_ (.CLK(clknet_4_4_0_clk),
    .D(net239),
    .RESET_B(_0018_),
    .Q(net41));
 sky130_fd_sc_hd__dfrtp_1 _1250_ (.CLK(clknet_4_0_0_clk),
    .D(net215),
    .RESET_B(_0019_),
    .Q(net42));
 sky130_fd_sc_hd__dfrtp_1 _1251_ (.CLK(clknet_4_5_0_clk),
    .D(_0206_),
    .RESET_B(_0020_),
    .Q(net43));
 sky130_fd_sc_hd__dfrtp_2 _1252_ (.CLK(clknet_4_2_0_clk),
    .D(net176),
    .RESET_B(_0021_),
    .Q(net44));
 sky130_fd_sc_hd__dfrtp_1 _1253_ (.CLK(clknet_4_4_0_clk),
    .D(_0208_),
    .RESET_B(_0022_),
    .Q(net55));
 sky130_fd_sc_hd__dfrtp_1 _1254_ (.CLK(clknet_4_4_0_clk),
    .D(net318),
    .RESET_B(_0023_),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_1 _1255_ (.CLK(clknet_4_0_0_clk),
    .D(net376),
    .RESET_B(_0024_),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _1256_ (.CLK(clknet_4_3_0_clk),
    .D(net339),
    .RESET_B(_0025_),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_2 _1257_ (.CLK(clknet_4_7_0_clk),
    .D(_0212_),
    .RESET_B(_0026_),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_2 _1258_ (.CLK(clknet_4_13_0_clk),
    .D(net161),
    .RESET_B(_0027_),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _1259_ (.CLK(clknet_4_5_0_clk),
    .D(_0214_),
    .RESET_B(_0028_),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _1260_ (.CLK(clknet_4_5_0_clk),
    .D(_0215_),
    .RESET_B(_0029_),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _1261_ (.CLK(clknet_4_8_0_clk),
    .D(_0216_),
    .RESET_B(_0030_),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_1 _1262_ (.CLK(clknet_4_0_0_clk),
    .D(net117),
    .RESET_B(_0031_),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _1263_ (.CLK(clknet_4_10_0_clk),
    .D(net186),
    .RESET_B(_0032_),
    .Q(net56));
 sky130_fd_sc_hd__dfrtp_1 _1264_ (.CLK(clknet_4_1_0_clk),
    .D(net196),
    .RESET_B(_0033_),
    .Q(net57));
 sky130_fd_sc_hd__dfrtp_1 _1265_ (.CLK(clknet_4_4_0_clk),
    .D(_0220_),
    .RESET_B(_0034_),
    .Q(net58));
 sky130_fd_sc_hd__dfrtp_1 _1266_ (.CLK(clknet_4_5_0_clk),
    .D(net291),
    .RESET_B(_0035_),
    .Q(net59));
 sky130_fd_sc_hd__dfrtp_1 _1267_ (.CLK(clknet_4_2_0_clk),
    .D(_0222_),
    .RESET_B(_0036_),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_1 _1268_ (.CLK(clknet_4_0_0_clk),
    .D(_0223_),
    .RESET_B(_0037_),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_1 _1269_ (.CLK(clknet_4_3_0_clk),
    .D(net127),
    .RESET_B(_0038_),
    .Q(net62));
 sky130_fd_sc_hd__dfrtp_1 _1270_ (.CLK(clknet_4_5_0_clk),
    .D(net255),
    .RESET_B(_0039_),
    .Q(net63));
 sky130_fd_sc_hd__dfrtp_1 _1271_ (.CLK(clknet_4_7_0_clk),
    .D(net251),
    .RESET_B(_0040_),
    .Q(net64));
 sky130_fd_sc_hd__dfrtp_2 _1272_ (.CLK(clknet_4_7_0_clk),
    .D(net272),
    .RESET_B(_0041_),
    .Q(net65));
 sky130_fd_sc_hd__dfrtp_2 _1273_ (.CLK(clknet_4_0_0_clk),
    .D(net119),
    .RESET_B(_0042_),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _1274_ (.CLK(clknet_4_0_0_clk),
    .D(net295),
    .RESET_B(_0043_),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_2 _1275_ (.CLK(clknet_4_7_0_clk),
    .D(net274),
    .RESET_B(_0044_),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_2 _1276_ (.CLK(clknet_4_7_0_clk),
    .D(net200),
    .RESET_B(_0045_),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _1277_ (.CLK(clknet_4_2_0_clk),
    .D(_0232_),
    .RESET_B(_0046_),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _1278_ (.CLK(clknet_4_13_0_clk),
    .D(_0233_),
    .RESET_B(_0047_),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _1279_ (.CLK(clknet_4_10_0_clk),
    .D(_0234_),
    .RESET_B(_0048_),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _1280_ (.CLK(clknet_4_5_0_clk),
    .D(_0235_),
    .RESET_B(_0049_),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _1281_ (.CLK(clknet_4_11_0_clk),
    .D(_0236_),
    .RESET_B(_0050_),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _1282_ (.CLK(clknet_4_0_0_clk),
    .D(_0237_),
    .RESET_B(_0051_),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _1283_ (.CLK(clknet_4_1_0_clk),
    .D(_0238_),
    .RESET_B(_0052_),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_1 _1284_ (.CLK(clknet_4_14_0_clk),
    .D(_0239_),
    .RESET_B(_0053_),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_1 _1285_ (.CLK(clknet_4_3_0_clk),
    .D(net387),
    .RESET_B(_0054_),
    .Q(\uart_tx_inst.i_data_valid ));
 sky130_fd_sc_hd__dfrtp_1 _1286_ (.CLK(clknet_4_9_0_clk),
    .D(net139),
    .RESET_B(_0055_),
    .Q(\uart_tx_inst.i_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1287_ (.CLK(clknet_4_8_0_clk),
    .D(net137),
    .RESET_B(_0056_),
    .Q(\uart_tx_inst.i_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1288_ (.CLK(clknet_4_3_0_clk),
    .D(net213),
    .RESET_B(_0057_),
    .Q(\uart_tx_inst.i_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1289_ (.CLK(clknet_4_3_0_clk),
    .D(net125),
    .RESET_B(_0058_),
    .Q(\uart_tx_inst.i_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1290_ (.CLK(clknet_4_9_0_clk),
    .D(net129),
    .RESET_B(_0059_),
    .Q(\uart_tx_inst.i_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1291_ (.CLK(clknet_4_3_0_clk),
    .D(net141),
    .RESET_B(_0060_),
    .Q(\uart_tx_inst.i_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1292_ (.CLK(clknet_4_2_0_clk),
    .D(net121),
    .RESET_B(_0061_),
    .Q(\uart_tx_inst.i_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1293_ (.CLK(clknet_4_8_0_clk),
    .D(net131),
    .RESET_B(_0062_),
    .Q(\uart_tx_inst.i_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1294_ (.CLK(clknet_4_6_0_clk),
    .D(net293),
    .RESET_B(_0063_),
    .Q(\cmd_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1295_ (.CLK(clknet_4_4_0_clk),
    .D(_0250_),
    .RESET_B(_0064_),
    .Q(\cmd_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1296_ (.CLK(clknet_4_4_0_clk),
    .D(_0251_),
    .RESET_B(_0065_),
    .Q(\cmd_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1297_ (.CLK(clknet_4_4_0_clk),
    .D(_0252_),
    .RESET_B(_0066_),
    .Q(\cmd_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1298_ (.CLK(clknet_4_4_0_clk),
    .D(_0253_),
    .RESET_B(_0067_),
    .Q(\cmd_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1299_ (.CLK(clknet_4_1_0_clk),
    .D(_0254_),
    .RESET_B(_0068_),
    .Q(\cmd_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1300_ (.CLK(clknet_4_1_0_clk),
    .D(_0255_),
    .RESET_B(_0069_),
    .Q(\cmd_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1301_ (.CLK(clknet_4_1_0_clk),
    .D(_0256_),
    .RESET_B(_0070_),
    .Q(\cmd_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1302_ (.CLK(clknet_4_6_0_clk),
    .D(net209),
    .RESET_B(_0071_),
    .Q(\addr_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1303_ (.CLK(clknet_4_5_0_clk),
    .D(_0258_),
    .RESET_B(_0072_),
    .Q(\addr_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1304_ (.CLK(clknet_4_5_0_clk),
    .D(net245),
    .RESET_B(_0073_),
    .Q(\addr_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1305_ (.CLK(clknet_4_6_0_clk),
    .D(net217),
    .RESET_B(_0074_),
    .Q(\addr_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1306_ (.CLK(clknet_4_1_0_clk),
    .D(net190),
    .RESET_B(_0075_),
    .Q(\addr_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1307_ (.CLK(clknet_4_7_0_clk),
    .D(net249),
    .RESET_B(_0076_),
    .Q(\addr_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1308_ (.CLK(clknet_4_5_0_clk),
    .D(net270),
    .RESET_B(_0077_),
    .Q(\addr_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1309_ (.CLK(clknet_4_4_0_clk),
    .D(_0264_),
    .RESET_B(_0078_),
    .Q(\addr_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1310_ (.CLK(clknet_4_7_0_clk),
    .D(_0265_),
    .RESET_B(_0079_),
    .Q(\addr_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1311_ (.CLK(clknet_4_9_0_clk),
    .D(net168),
    .RESET_B(_0080_),
    .Q(\addr_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1312_ (.CLK(clknet_4_7_0_clk),
    .D(net232),
    .RESET_B(_0081_),
    .Q(\addr_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1313_ (.CLK(clknet_4_9_0_clk),
    .D(net166),
    .RESET_B(_0082_),
    .Q(\addr_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1314_ (.CLK(clknet_4_4_0_clk),
    .D(net230),
    .RESET_B(_0083_),
    .Q(\addr_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1315_ (.CLK(clknet_4_0_0_clk),
    .D(net188),
    .RESET_B(_0084_),
    .Q(\addr_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1316_ (.CLK(clknet_4_5_0_clk),
    .D(net260),
    .RESET_B(_0085_),
    .Q(\addr_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1317_ (.CLK(clknet_4_0_0_clk),
    .D(net180),
    .RESET_B(_0086_),
    .Q(\addr_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1318_ (.CLK(clknet_4_4_0_clk),
    .D(net234),
    .RESET_B(_0087_),
    .Q(\data_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1319_ (.CLK(clknet_4_5_0_clk),
    .D(_0274_),
    .RESET_B(_0088_),
    .Q(\data_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1320_ (.CLK(clknet_4_4_0_clk),
    .D(_0275_),
    .RESET_B(_0089_),
    .Q(\data_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1321_ (.CLK(clknet_4_6_0_clk),
    .D(_0276_),
    .RESET_B(_0090_),
    .Q(\data_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1322_ (.CLK(clknet_4_5_0_clk),
    .D(net308),
    .RESET_B(_0091_),
    .Q(\data_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1323_ (.CLK(clknet_4_7_0_clk),
    .D(_0278_),
    .RESET_B(_0092_),
    .Q(\data_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1324_ (.CLK(clknet_4_5_0_clk),
    .D(net298),
    .RESET_B(_0093_),
    .Q(\data_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1325_ (.CLK(clknet_4_5_0_clk),
    .D(net262),
    .RESET_B(_0094_),
    .Q(\data_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1326_ (.CLK(clknet_4_8_0_clk),
    .D(net253),
    .RESET_B(_0095_),
    .Q(\data_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1327_ (.CLK(clknet_4_1_0_clk),
    .D(net170),
    .RESET_B(_0096_),
    .Q(\data_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1328_ (.CLK(clknet_4_8_0_clk),
    .D(net287),
    .RESET_B(_0097_),
    .Q(\data_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1329_ (.CLK(clknet_4_1_0_clk),
    .D(net153),
    .RESET_B(_0098_),
    .Q(\data_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1330_ (.CLK(clknet_4_4_0_clk),
    .D(net243),
    .RESET_B(_0099_),
    .Q(\data_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1331_ (.CLK(clknet_4_4_0_clk),
    .D(_0286_),
    .RESET_B(_0100_),
    .Q(\data_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1332_ (.CLK(clknet_4_2_0_clk),
    .D(net178),
    .RESET_B(_0101_),
    .Q(\data_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1333_ (.CLK(clknet_4_0_0_clk),
    .D(net219),
    .RESET_B(_0102_),
    .Q(\data_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1334_ (.CLK(clknet_4_2_0_clk),
    .D(_0289_),
    .RESET_B(_0103_),
    .Q(\data_reg[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1335_ (.CLK(clknet_4_5_0_clk),
    .D(_0290_),
    .RESET_B(_0104_),
    .Q(\data_reg[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1336_ (.CLK(clknet_4_7_0_clk),
    .D(net258),
    .RESET_B(_0105_),
    .Q(\data_reg[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1337_ (.CLK(clknet_4_7_0_clk),
    .D(_0292_),
    .RESET_B(_0106_),
    .Q(\data_reg[19] ));
 sky130_fd_sc_hd__dfrtp_1 _1338_ (.CLK(clknet_4_1_0_clk),
    .D(_0293_),
    .RESET_B(_0107_),
    .Q(\data_reg[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1339_ (.CLK(clknet_4_0_0_clk),
    .D(_0294_),
    .RESET_B(_0108_),
    .Q(\data_reg[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1340_ (.CLK(clknet_4_5_0_clk),
    .D(_0295_),
    .RESET_B(_0109_),
    .Q(\data_reg[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1341_ (.CLK(clknet_4_7_0_clk),
    .D(net207),
    .RESET_B(_0110_),
    .Q(\data_reg[23] ));
 sky130_fd_sc_hd__dfrtp_4 _1342_ (.CLK(clknet_4_3_0_clk),
    .D(_0297_),
    .RESET_B(_0111_),
    .Q(\byte_count[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1343_ (.CLK(clknet_4_3_0_clk),
    .D(_0298_),
    .RESET_B(_0112_),
    .Q(\byte_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1344_ (.CLK(clknet_4_3_0_clk),
    .D(_0299_),
    .RESET_B(_0113_),
    .Q(\byte_count[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1345_ (.CLK(clknet_4_3_0_clk),
    .D(_0300_),
    .RESET_B(_0114_),
    .Q(\byte_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1346_ (.CLK(clknet_4_6_0_clk),
    .D(_0301_),
    .RESET_B(_0115_),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1347_ (.CLK(clknet_4_6_0_clk),
    .D(_0302_),
    .RESET_B(_0116_),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1348_ (.CLK(clknet_4_6_0_clk),
    .D(_0303_),
    .RESET_B(_0117_),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfstp_1 _1349_ (.CLK(clknet_4_11_0_clk),
    .D(net2),
    .SET_B(_0118_),
    .Q(\uart_rx_inst.rx_sync_1 ));
 sky130_fd_sc_hd__dfrtp_1 _1350_ (.CLK(clknet_4_15_0_clk),
    .D(_0001_),
    .RESET_B(_0119_),
    .Q(\uart_rx_inst.receiving ));
 sky130_fd_sc_hd__dfrtp_1 _1351_ (.CLK(clknet_4_13_0_clk),
    .D(_0304_),
    .RESET_B(_0120_),
    .Q(\uart_rx_inst.clock_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1352_ (.CLK(clknet_4_13_0_clk),
    .D(net349),
    .RESET_B(_0121_),
    .Q(\uart_rx_inst.clock_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1353_ (.CLK(clknet_4_13_0_clk),
    .D(net341),
    .RESET_B(_0122_),
    .Q(\uart_rx_inst.clock_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1354_ (.CLK(clknet_4_13_0_clk),
    .D(net327),
    .RESET_B(_0123_),
    .Q(\uart_rx_inst.clock_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1355_ (.CLK(clknet_4_15_0_clk),
    .D(net381),
    .RESET_B(_0124_),
    .Q(\uart_rx_inst.clock_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1356_ (.CLK(clknet_4_15_0_clk),
    .D(net337),
    .RESET_B(_0125_),
    .Q(\uart_rx_inst.clock_count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1357_ (.CLK(clknet_4_15_0_clk),
    .D(_0310_),
    .RESET_B(_0126_),
    .Q(\uart_rx_inst.clock_count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1358_ (.CLK(clknet_4_15_0_clk),
    .D(net329),
    .RESET_B(_0127_),
    .Q(\uart_rx_inst.clock_count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1359_ (.CLK(clknet_4_15_0_clk),
    .D(_0312_),
    .RESET_B(_0128_),
    .Q(\uart_rx_inst.clock_count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1360_ (.CLK(clknet_4_15_0_clk),
    .D(net310),
    .RESET_B(_0129_),
    .Q(\uart_rx_inst.clock_count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1361_ (.CLK(clknet_4_15_0_clk),
    .D(net358),
    .RESET_B(_0130_),
    .Q(\uart_rx_inst.clock_count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1362_ (.CLK(clknet_4_15_0_clk),
    .D(net314),
    .RESET_B(_0131_),
    .Q(\uart_rx_inst.clock_count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1363_ (.CLK(clknet_4_15_0_clk),
    .D(_0316_),
    .RESET_B(_0132_),
    .Q(\uart_rx_inst.clock_count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1364_ (.CLK(clknet_4_13_0_clk),
    .D(net325),
    .RESET_B(_0133_),
    .Q(\uart_rx_inst.clock_count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1365_ (.CLK(clknet_4_13_0_clk),
    .D(net346),
    .RESET_B(_0134_),
    .Q(\uart_rx_inst.clock_count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1366_ (.CLK(clknet_4_13_0_clk),
    .D(_0319_),
    .RESET_B(_0135_),
    .Q(\uart_rx_inst.clock_count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1367_ (.CLK(clknet_4_15_0_clk),
    .D(_0320_),
    .RESET_B(_0136_),
    .Q(\uart_rx_inst.bit_index[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1368_ (.CLK(clknet_4_14_0_clk),
    .D(_0321_),
    .RESET_B(_0137_),
    .Q(\uart_rx_inst.bit_index[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1369_ (.CLK(clknet_4_15_0_clk),
    .D(_0322_),
    .RESET_B(_0138_),
    .Q(\uart_rx_inst.bit_index[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1370_ (.CLK(clknet_4_12_0_clk),
    .D(net194),
    .RESET_B(_0139_),
    .Q(\uart_rx_inst.bit_index[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1371_ (.CLK(clknet_4_12_0_clk),
    .D(net149),
    .RESET_B(_0140_),
    .Q(\uart_rx_inst.o_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1372_ (.CLK(clknet_4_12_0_clk),
    .D(net133),
    .RESET_B(_0141_),
    .Q(\uart_rx_inst.o_data[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1373_ (.CLK(clknet_4_14_0_clk),
    .D(net184),
    .RESET_B(_0142_),
    .Q(\uart_rx_inst.o_data[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1374_ (.CLK(clknet_4_12_0_clk),
    .D(net267),
    .RESET_B(_0143_),
    .Q(\uart_rx_inst.o_data[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1375_ (.CLK(clknet_4_14_0_clk),
    .D(net223),
    .RESET_B(_0144_),
    .Q(\uart_rx_inst.o_data[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1376_ (.CLK(clknet_4_12_0_clk),
    .D(net151),
    .RESET_B(_0145_),
    .Q(\uart_rx_inst.o_data[5] ));
 sky130_fd_sc_hd__dfrtp_4 _1377_ (.CLK(clknet_4_12_0_clk),
    .D(net145),
    .RESET_B(_0146_),
    .Q(\uart_rx_inst.o_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1378_ (.CLK(clknet_4_14_0_clk),
    .D(net182),
    .RESET_B(_0147_),
    .Q(\uart_rx_inst.o_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1379_ (.CLK(clknet_4_12_0_clk),
    .D(_0000_),
    .RESET_B(_0148_),
    .Q(\uart_rx_inst.o_data_valid ));
 sky130_fd_sc_hd__dfrtp_1 _1380_ (.CLK(clknet_4_9_0_clk),
    .D(net241),
    .RESET_B(_0149_),
    .Q(\uart_tx_inst.shift_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1381_ (.CLK(clknet_4_8_0_clk),
    .D(net159),
    .RESET_B(_0150_),
    .Q(\uart_tx_inst.shift_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1382_ (.CLK(clknet_4_8_0_clk),
    .D(net135),
    .RESET_B(_0151_),
    .Q(\uart_tx_inst.shift_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1383_ (.CLK(clknet_4_3_0_clk),
    .D(net221),
    .RESET_B(_0152_),
    .Q(\uart_tx_inst.shift_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1384_ (.CLK(clknet_4_9_0_clk),
    .D(net202),
    .RESET_B(_0153_),
    .Q(\uart_tx_inst.shift_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1385_ (.CLK(clknet_4_2_0_clk),
    .D(net157),
    .RESET_B(_0154_),
    .Q(\uart_tx_inst.shift_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1386_ (.CLK(clknet_4_2_0_clk),
    .D(net155),
    .RESET_B(_0155_),
    .Q(\uart_tx_inst.shift_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1387_ (.CLK(clknet_4_8_0_clk),
    .D(net143),
    .RESET_B(_0156_),
    .Q(\uart_tx_inst.shift_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1388_ (.CLK(clknet_4_8_0_clk),
    .D(net123),
    .RESET_B(_0157_),
    .Q(\uart_tx_inst.shift_reg[9] ));
 sky130_fd_sc_hd__dfstp_1 _1389_ (.CLK(clknet_4_14_0_clk),
    .D(net115),
    .SET_B(_0158_),
    .Q(\uart_rx_inst.rx_sync_2 ));
 sky130_fd_sc_hd__dfrtp_1 _1390_ (.CLK(clknet_4_9_0_clk),
    .D(_0002_),
    .RESET_B(_0159_),
    .Q(\uart_tx_inst.transmitting ));
 sky130_fd_sc_hd__dfstp_1 _1391_ (.CLK(clknet_4_10_0_clk),
    .D(net420),
    .SET_B(_0160_),
    .Q(net37));
 sky130_fd_sc_hd__dfrtp_1 _1392_ (.CLK(clknet_4_11_0_clk),
    .D(net395),
    .RESET_B(_0161_),
    .Q(\uart_tx_inst.clock_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1393_ (.CLK(clknet_4_11_0_clk),
    .D(net383),
    .RESET_B(_0162_),
    .Q(\uart_tx_inst.clock_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1394_ (.CLK(clknet_4_11_0_clk),
    .D(net363),
    .RESET_B(_0163_),
    .Q(\uart_tx_inst.clock_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1395_ (.CLK(clknet_4_11_0_clk),
    .D(net316),
    .RESET_B(_0164_),
    .Q(\uart_tx_inst.clock_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1396_ (.CLK(clknet_4_10_0_clk),
    .D(net369),
    .RESET_B(_0165_),
    .Q(\uart_tx_inst.clock_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1397_ (.CLK(clknet_4_10_0_clk),
    .D(net409),
    .RESET_B(_0166_),
    .Q(\uart_tx_inst.clock_count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1398_ (.CLK(clknet_4_10_0_clk),
    .D(net360),
    .RESET_B(_0167_),
    .Q(\uart_tx_inst.clock_count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1399_ (.CLK(clknet_4_10_0_clk),
    .D(net393),
    .RESET_B(_0168_),
    .Q(\uart_tx_inst.clock_count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1400_ (.CLK(clknet_4_10_0_clk),
    .D(net403),
    .RESET_B(_0169_),
    .Q(\uart_tx_inst.clock_count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1401_ (.CLK(clknet_4_10_0_clk),
    .D(net398),
    .RESET_B(_0170_),
    .Q(\uart_tx_inst.clock_count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1402_ (.CLK(clknet_4_10_0_clk),
    .D(net367),
    .RESET_B(_0171_),
    .Q(\uart_tx_inst.clock_count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1403_ (.CLK(clknet_4_10_0_clk),
    .D(net401),
    .RESET_B(_0172_),
    .Q(\uart_tx_inst.clock_count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1404_ (.CLK(clknet_4_10_0_clk),
    .D(net332),
    .RESET_B(_0173_),
    .Q(\uart_tx_inst.clock_count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1405_ (.CLK(clknet_4_11_0_clk),
    .D(net406),
    .RESET_B(_0174_),
    .Q(\uart_tx_inst.clock_count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1406_ (.CLK(clknet_4_11_0_clk),
    .D(net334),
    .RESET_B(_0175_),
    .Q(\uart_tx_inst.clock_count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1407_ (.CLK(clknet_4_11_0_clk),
    .D(net303),
    .RESET_B(_0176_),
    .Q(\uart_tx_inst.clock_count[15] ));
 sky130_fd_sc_hd__dfrtp_2 _1408_ (.CLK(clknet_4_8_0_clk),
    .D(_0358_),
    .RESET_B(_0177_),
    .Q(\uart_tx_inst.bit_index[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1409_ (.CLK(clknet_4_8_0_clk),
    .D(net385),
    .RESET_B(_0178_),
    .Q(\uart_tx_inst.bit_index[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1410_ (.CLK(clknet_4_8_0_clk),
    .D(net378),
    .RESET_B(_0179_),
    .Q(\uart_tx_inst.bit_index[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1411_ (.CLK(clknet_4_8_0_clk),
    .D(net389),
    .RESET_B(_0180_),
    .Q(\uart_tx_inst.bit_index[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1412_ (.CLK(clknet_4_12_0_clk),
    .D(net164),
    .RESET_B(_0181_),
    .Q(\uart_rx_inst.shift_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1413_ (.CLK(clknet_4_14_0_clk),
    .D(_0363_),
    .RESET_B(_0182_),
    .Q(\uart_rx_inst.shift_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1414_ (.CLK(clknet_4_14_0_clk),
    .D(net344),
    .RESET_B(_0183_),
    .Q(\uart_rx_inst.shift_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1415_ (.CLK(clknet_4_12_0_clk),
    .D(_0365_),
    .RESET_B(_0184_),
    .Q(\uart_rx_inst.shift_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1416_ (.CLK(clknet_4_14_0_clk),
    .D(_0366_),
    .RESET_B(_0185_),
    .Q(\uart_rx_inst.shift_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1417_ (.CLK(clknet_4_12_0_clk),
    .D(net174),
    .RESET_B(_0186_),
    .Q(\uart_rx_inst.shift_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1418_ (.CLK(clknet_4_13_0_clk),
    .D(net227),
    .RESET_B(_0187_),
    .Q(\uart_rx_inst.shift_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1419_ (.CLK(clknet_4_14_0_clk),
    .D(_0369_),
    .RESET_B(_0188_),
    .Q(\uart_rx_inst.shift_reg[7] ));
 sky130_fd_sc_hd__buf_1 _1420_ (.A(net54),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__buf_8 fanout100 (.A(net106),
    .X(net100));
 sky130_fd_sc_hd__buf_8 fanout101 (.A(net106),
    .X(net101));
 sky130_fd_sc_hd__buf_8 fanout102 (.A(net106),
    .X(net102));
 sky130_fd_sc_hd__buf_4 fanout103 (.A(net106),
    .X(net103));
 sky130_fd_sc_hd__buf_8 fanout104 (.A(net106),
    .X(net104));
 sky130_fd_sc_hd__buf_4 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_8 fanout106 (.A(net3),
    .X(net106));
 sky130_fd_sc_hd__buf_6 fanout107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__buf_4 fanout108 (.A(net3),
    .X(net108));
 sky130_fd_sc_hd__buf_8 fanout109 (.A(net3),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_8 fanout110 (.A(net3),
    .X(net110));
 sky130_fd_sc_hd__buf_8 fanout111 (.A(net114),
    .X(net111));
 sky130_fd_sc_hd__buf_8 fanout112 (.A(net114),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__buf_4 fanout114 (.A(net3),
    .X(net114));
 sky130_fd_sc_hd__buf_6 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__buf_6 fanout90 (.A(_0612_),
    .X(net90));
 sky130_fd_sc_hd__buf_4 fanout91 (.A(net92),
    .X(net91));
 sky130_fd_sc_hd__buf_4 fanout92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_8 fanout93 (.A(_0572_),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_8 fanout96 (.A(net414),
    .X(net96));
 sky130_fd_sc_hd__buf_4 fanout97 (.A(net355),
    .X(net97));
 sky130_fd_sc_hd__buf_2 fanout98 (.A(net355),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_8 fanout99 (.A(net205),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net424),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\uart_tx_inst.i_data[3] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net42),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_0205_),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\addr_reg[3] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_0260_),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\data_reg[15] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0288_),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\uart_tx_inst.shift_reg[4] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0335_),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\uart_rx_inst.shift_reg[4] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0328_),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0244_),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net60),
    .X(net224));
 sky130_fd_sc_hd__buf_2 hold111 (.A(net433),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0406_),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_0368_),
    .X(net227));
 sky130_fd_sc_hd__buf_2 hold114 (.A(net430),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\addr_reg[12] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_0269_),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\addr_reg[10] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_0267_),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\data_reg[0] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\data_reg[16] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0273_),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net48),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(net38),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0192_),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(net41),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_0204_),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\uart_tx_inst.shift_reg[1] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_0332_),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\data_reg[12] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0285_),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0224_),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\addr_reg[2] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_0259_),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(net61),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 hold133 (.A(\uart_rx_inst.o_data_valid ),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 hold134 (.A(_0530_),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0262_),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\data_reg[18] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0226_),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\data_reg[8] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_0281_),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\uart_tx_inst.i_data[4] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\data_reg[17] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_0225_),
    .X(net255));
 sky130_fd_sc_hd__buf_2 hold142 (.A(\byte_count[3] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_0577_),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_0291_),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\addr_reg[14] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0271_),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\data_reg[7] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0280_),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 hold149 (.A(net432),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0245_),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_0583_),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(net39),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\uart_rx_inst.shift_reg[3] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_0327_),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(net46),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\addr_reg[6] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_0263_),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\data_reg[19] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0227_),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\data_reg[22] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\uart_tx_inst.i_data[7] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_0230_),
    .X(net274));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold161 (.A(\byte_count[1] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(net55),
    .X(net276));
 sky130_fd_sc_hd__buf_1 hold163 (.A(\uart_rx_inst.o_data[3] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(net43),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(net58),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\addr_reg[7] ),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_2 hold167 (.A(\uart_rx_inst.o_data[6] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(net47),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(net85),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0248_),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(net84),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\cmd_reg[5] ),
    .X(net285));
 sky130_fd_sc_hd__buf_2 hold172 (.A(\uart_rx_inst.o_data[2] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_0283_),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_2 hold174 (.A(\uart_rx_inst.o_data[4] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(net50),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\data_reg[13] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_0221_),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\cmd_reg[0] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_0249_),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\uart_rx_inst.shift_reg[1] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\data_reg[21] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_0229_),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(net51),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\data_reg[6] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_0279_),
    .X(net298));
 sky130_fd_sc_hd__buf_2 hold185 (.A(\state[0] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_0536_),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\cmd_reg[7] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\uart_tx_inst.clock_count[15] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_0357_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0325_),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\cmd_reg[2] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\cmd_reg[4] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\cmd_reg[6] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\data_reg[4] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_0277_),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\uart_rx_inst.clock_count[9] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_0313_),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\cmd_reg[3] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(net83),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\uart_rx_inst.clock_count[11] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\data_reg[9] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\uart_tx_inst.i_data[2] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_0315_),
    .X(net314));
 sky130_fd_sc_hd__buf_1 hold201 (.A(\uart_tx_inst.clock_count[3] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_0345_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\data_reg[1] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_0209_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(net81),
    .X(net319));
 sky130_fd_sc_hd__buf_2 hold206 (.A(\state[2] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_0532_),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_0569_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\cmd_reg[1] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0334_),
    .X(net135));
 sky130_fd_sc_hd__buf_1 hold210 (.A(\uart_rx_inst.clock_count[13] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_0317_),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\uart_rx_inst.clock_count[3] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_0307_),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\uart_rx_inst.clock_count[7] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_0311_),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\addr_reg[1] ),
    .X(net330));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold217 (.A(\uart_tx_inst.clock_count[12] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_0354_),
    .X(net332));
 sky130_fd_sc_hd__buf_1 hold219 (.A(\uart_tx_inst.clock_count[14] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\uart_tx_inst.i_data[1] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_0356_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(net45),
    .X(net335));
 sky130_fd_sc_hd__buf_1 hold222 (.A(\uart_rx_inst.clock_count[5] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_0309_),
    .X(net337));
 sky130_fd_sc_hd__buf_1 hold224 (.A(net429),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0211_),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\uart_rx_inst.clock_count[2] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_0306_),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\byte_count[1] ),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_4 hold229 (.A(net426),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_0242_),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_0364_),
    .X(net344));
 sky130_fd_sc_hd__buf_1 hold231 (.A(\uart_rx_inst.clock_count[14] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0318_),
    .X(net346));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold233 (.A(\uart_rx_inst.clock_count[1] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_0517_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_0305_),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\uart_rx_inst.clock_count[15] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_0389_),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_0396_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_0397_),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\uart_tx_inst.i_data[0] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0414_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\uart_rx_inst.receiving ),
    .X(net355));
 sky130_fd_sc_hd__buf_2 hold242 (.A(net435),
    .X(net356));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold243 (.A(\uart_rx_inst.clock_count[10] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_0314_),
    .X(net358));
 sky130_fd_sc_hd__buf_1 hold245 (.A(\uart_tx_inst.clock_count[6] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_0348_),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(net79),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\uart_tx_inst.clock_count[2] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_0344_),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0241_),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(net72),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(net75),
    .X(net365));
 sky130_fd_sc_hd__buf_1 hold252 (.A(\uart_tx_inst.clock_count[10] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_0352_),
    .X(net367));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold254 (.A(\uart_tx_inst.clock_count[4] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_0346_),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(net78),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(net88),
    .X(net371));
 sky130_fd_sc_hd__buf_1 hold258 (.A(net428),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(net73),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\uart_tx_inst.i_data[5] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(net76),
    .X(net374));
 sky130_fd_sc_hd__buf_1 hold261 (.A(net434),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_0210_),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_2 hold263 (.A(\uart_tx_inst.bit_index[2] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_0360_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(net71),
    .X(net379));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold266 (.A(\uart_rx_inst.clock_count[4] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_0308_),
    .X(net381));
 sky130_fd_sc_hd__buf_1 hold268 (.A(\uart_tx_inst.clock_count[1] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_0343_),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0246_),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 hold270 (.A(\uart_tx_inst.bit_index[1] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(_0359_),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_2 hold272 (.A(net437),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_0240_),
    .X(net387));
 sky130_fd_sc_hd__buf_1 hold274 (.A(\uart_tx_inst.bit_index[3] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_0361_),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(net74),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\uart_tx_inst.clock_count[7] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_0461_),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(_0349_),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\uart_tx_inst.shift_reg[8] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\uart_tx_inst.clock_count[0] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_0342_),
    .X(net395));
 sky130_fd_sc_hd__buf_1 hold282 (.A(\uart_tx_inst.clock_count[9] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_0458_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_0351_),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\uart_rx_inst.clock_count[0] ),
    .X(net399));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold286 (.A(\uart_tx_inst.clock_count[11] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_0353_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\uart_tx_inst.clock_count[8] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_0350_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_0339_),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\uart_tx_inst.clock_count[13] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_0449_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_0355_),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\uart_tx_inst.clock_count[5] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_0464_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_0347_),
    .X(net409));
 sky130_fd_sc_hd__buf_2 hold296 (.A(\uart_tx_inst.o_ready ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_0189_),
    .X(net411));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold298 (.A(\uart_rx_inst.clock_count[8] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_0390_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_0217_),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\uart_rx_inst.shift_reg[6] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\uart_tx_inst.transmitting ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\uart_rx_inst.clock_count[6] ),
    .X(net415));
 sky130_fd_sc_hd__buf_1 hold302 (.A(\uart_tx_inst.bit_index[0] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(net54),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\state[1] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(net37),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_0341_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\state[2] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\byte_count[3] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\state[0] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_0330_),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\uart_rx_inst.rx_sync_1 ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\uart_tx_inst.shift_reg[3] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\uart_rx_inst.bit_index[1] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\uart_rx_inst.bit_index[0] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\uart_rx_inst.clock_count[12] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\data_reg[3] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\uart_rx_inst.o_data[0] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\uart_rx_inst.o_data[7] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\uart_rx_inst.o_data[5] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\uart_rx_inst.bit_index[2] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\addr_reg[8] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\data_reg[2] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\state[1] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\uart_rx_inst.rx_sync_2 ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\uart_tx_inst.i_data_valid ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\uart_rx_inst.o_data[1] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_0200_),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\uart_rx_inst.shift_reg[0] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_0324_),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\uart_rx_inst.shift_reg[5] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_0329_),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\data_reg[11] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0284_),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\data_reg[20] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\uart_tx_inst.shift_reg[7] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0338_),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\uart_tx_inst.shift_reg[6] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_0337_),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\uart_tx_inst.shift_reg[2] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0333_),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\data_reg[5] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0213_),
    .X(net161));
 sky130_fd_sc_hd__buf_2 hold48 (.A(net436),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0402_),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_0228_),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0362_),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\addr_reg[11] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0268_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\addr_reg[9] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0266_),
    .X(net168));
 sky130_fd_sc_hd__buf_2 hold55 (.A(net438),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0282_),
    .X(net170));
 sky130_fd_sc_hd__buf_2 hold57 (.A(net427),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0408_),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0409_),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\uart_tx_inst.i_data[6] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0367_),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\addr_reg[15] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0207_),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\data_reg[14] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0287_),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_4 hold65 (.A(net431),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0272_),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\uart_rx_inst.shift_reg[7] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0331_),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\uart_rx_inst.shift_reg[2] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_0247_),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0326_),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\data_reg[10] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0218_),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\addr_reg[13] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0270_),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\addr_reg[4] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0261_),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\addr_reg[5] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0197_),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\uart_rx_inst.bit_index[3] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\uart_tx_inst.shift_reg[9] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0323_),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net57),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0219_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net40),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0203_),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\data_reg[23] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0231_),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\uart_tx_inst.shift_reg[5] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0336_),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net53),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0340_),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0201_),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_2 hold91 (.A(\byte_count[0] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0571_),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0296_),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\addr_reg[0] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_0257_),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 hold96 (.A(\byte_count[2] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0591_),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0603_),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0243_),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(i_start_rx),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(wb_dat_i[14]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(wb_dat_i[15]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(wb_dat_i[16]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(wb_dat_i[17]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(wb_dat_i[18]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(wb_dat_i[19]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(wb_dat_i[1]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(wb_dat_i[20]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(wb_dat_i[21]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(wb_dat_i[22]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(i_uart_rx),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(wb_dat_i[23]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(wb_dat_i[24]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(wb_dat_i[25]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(wb_dat_i[26]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(wb_dat_i[27]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(wb_dat_i[28]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(wb_dat_i[29]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(wb_dat_i[2]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(wb_dat_i[30]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(wb_dat_i[31]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(rst),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(wb_dat_i[3]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(wb_dat_i[4]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(wb_dat_i[5]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(wb_dat_i[6]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(wb_dat_i[7]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(wb_dat_i[8]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(wb_dat_i[9]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input4 (.A(wb_ack_i),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(wb_dat_i[0]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(wb_dat_i[10]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(wb_dat_i[11]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(wb_dat_i[12]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(wb_dat_i[13]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 max_cap95 (.A(_0392_),
    .X(net95));
 sky130_fd_sc_hd__buf_12 output37 (.A(net37),
    .X(o_uart_tx));
 sky130_fd_sc_hd__buf_12 output38 (.A(net38),
    .X(wb_adr_o[0]));
 sky130_fd_sc_hd__buf_12 output39 (.A(net39),
    .X(wb_adr_o[10]));
 sky130_fd_sc_hd__buf_12 output40 (.A(net40),
    .X(wb_adr_o[11]));
 sky130_fd_sc_hd__buf_12 output41 (.A(net41),
    .X(wb_adr_o[12]));
 sky130_fd_sc_hd__buf_12 output42 (.A(net42),
    .X(wb_adr_o[13]));
 sky130_fd_sc_hd__buf_12 output43 (.A(net43),
    .X(wb_adr_o[14]));
 sky130_fd_sc_hd__buf_12 output44 (.A(net44),
    .X(wb_adr_o[15]));
 sky130_fd_sc_hd__buf_12 output45 (.A(net45),
    .X(wb_adr_o[1]));
 sky130_fd_sc_hd__buf_12 output46 (.A(net46),
    .X(wb_adr_o[2]));
 sky130_fd_sc_hd__buf_12 output47 (.A(net47),
    .X(wb_adr_o[3]));
 sky130_fd_sc_hd__buf_12 output48 (.A(net48),
    .X(wb_adr_o[4]));
 sky130_fd_sc_hd__buf_12 output49 (.A(net49),
    .X(wb_adr_o[5]));
 sky130_fd_sc_hd__buf_12 output50 (.A(net50),
    .X(wb_adr_o[6]));
 sky130_fd_sc_hd__buf_12 output51 (.A(net51),
    .X(wb_adr_o[7]));
 sky130_fd_sc_hd__buf_12 output52 (.A(net52),
    .X(wb_adr_o[8]));
 sky130_fd_sc_hd__buf_12 output53 (.A(net53),
    .X(wb_adr_o[9]));
 sky130_fd_sc_hd__buf_12 output54 (.A(net54),
    .X(wb_cyc_o));
 sky130_fd_sc_hd__buf_12 output55 (.A(net55),
    .X(wb_dat_o[0]));
 sky130_fd_sc_hd__buf_12 output56 (.A(net56),
    .X(wb_dat_o[10]));
 sky130_fd_sc_hd__buf_12 output57 (.A(net57),
    .X(wb_dat_o[11]));
 sky130_fd_sc_hd__buf_12 output58 (.A(net58),
    .X(wb_dat_o[12]));
 sky130_fd_sc_hd__buf_12 output59 (.A(net59),
    .X(wb_dat_o[13]));
 sky130_fd_sc_hd__buf_12 output60 (.A(net60),
    .X(wb_dat_o[14]));
 sky130_fd_sc_hd__buf_12 output61 (.A(net61),
    .X(wb_dat_o[15]));
 sky130_fd_sc_hd__buf_12 output62 (.A(net62),
    .X(wb_dat_o[16]));
 sky130_fd_sc_hd__buf_12 output63 (.A(net63),
    .X(wb_dat_o[17]));
 sky130_fd_sc_hd__buf_12 output64 (.A(net64),
    .X(wb_dat_o[18]));
 sky130_fd_sc_hd__buf_12 output65 (.A(net65),
    .X(wb_dat_o[19]));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(wb_dat_o[1]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(wb_dat_o[20]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(wb_dat_o[21]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(wb_dat_o[22]));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(wb_dat_o[23]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(wb_dat_o[24]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net72),
    .X(wb_dat_o[25]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(wb_dat_o[26]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(wb_dat_o[27]));
 sky130_fd_sc_hd__buf_12 output75 (.A(net75),
    .X(wb_dat_o[28]));
 sky130_fd_sc_hd__buf_12 output76 (.A(net76),
    .X(wb_dat_o[29]));
 sky130_fd_sc_hd__buf_12 output77 (.A(net77),
    .X(wb_dat_o[2]));
 sky130_fd_sc_hd__buf_12 output78 (.A(net78),
    .X(wb_dat_o[30]));
 sky130_fd_sc_hd__buf_12 output79 (.A(net79),
    .X(wb_dat_o[31]));
 sky130_fd_sc_hd__buf_12 output80 (.A(net80),
    .X(wb_dat_o[3]));
 sky130_fd_sc_hd__buf_12 output81 (.A(net81),
    .X(wb_dat_o[4]));
 sky130_fd_sc_hd__buf_12 output82 (.A(net82),
    .X(wb_dat_o[5]));
 sky130_fd_sc_hd__buf_12 output83 (.A(net83),
    .X(wb_dat_o[6]));
 sky130_fd_sc_hd__buf_12 output84 (.A(net84),
    .X(wb_dat_o[7]));
 sky130_fd_sc_hd__buf_12 output85 (.A(net85),
    .X(wb_dat_o[8]));
 sky130_fd_sc_hd__buf_12 output86 (.A(net86),
    .X(wb_dat_o[9]));
 sky130_fd_sc_hd__buf_12 output87 (.A(net87),
    .X(wb_stb_o));
 sky130_fd_sc_hd__buf_12 output88 (.A(net88),
    .X(wb_we_o));
 sky130_fd_sc_hd__buf_1 wire94 (.A(_0555_),
    .X(net94));
endmodule

